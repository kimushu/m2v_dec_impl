// demo_de0_sys.v

// Generated using ACDS version 11.1sp2 259 at 2012.08.24.21:44:24

`timescale 1 ps / 1 ps
module demo_de0_sys (
		input  wire        pll_areset_export,          //    pll_areset.export
		output wire [21:0] flash_tcm_address_out,      //         flash.tcm_address_out
		output wire        flash_tcm_read_n_out,       //              .tcm_read_n_out
		output wire        flash_tcm_write_n_out,      //              .tcm_write_n_out
		inout  wire [15:0] flash_tcm_data_out,         //              .tcm_data_out
		output wire        flash_tcm_chipselect_n_out, //              .tcm_chipselect_n_out
		output wire        pll_phasedone_export,       // pll_phasedone.export
		output wire [11:0] sdr_addr,                   //           sdr.addr
		output wire [1:0]  sdr_ba,                     //              .ba
		output wire        sdr_cas_n,                  //              .cas_n
		output wire        sdr_cke,                    //              .cke
		output wire        sdr_cs_n,                   //              .cs_n
		inout  wire [15:0] sdr_dq,                     //              .dq
		output wire [1:0]  sdr_dqm,                    //              .dqm
		output wire        sdr_ras_n,                  //              .ras_n
		output wire        sdr_we_n,                   //              .we_n
		output wire        sdrclk_clk,                 //        sdrclk.clk
		input  wire        reset_reset_n,              //         reset.reset_n
		output wire        lcd_reset_n,                //           lcd.reset_n
		output wire        lcd_cs,                     //              .cs
		output wire        lcd_rs,                     //              .rs
		inout  wire [15:0] lcd_data,                   //              .data
		output wire        lcd_write_n,                //              .write_n
		output wire        lcd_read_n,                 //              .read_n
		output wire [3:0]  hd_a,                       //            hd.a
		output wire [3:0]  hd_b,                       //              .b
		output wire [3:0]  hd_c,                       //              .c
		output wire [3:0]  hd_d,                       //              .d
		output wire [3:0]  hd_e,                       //              .e
		output wire [3:0]  hd_f,                       //              .f
		output wire [3:0]  hd_g,                       //              .g
		output wire [3:0]  hd_dp,                      //              .dp
		input  wire        clk_clk,                    //           clk.clk
		output wire        pll_locked_export,          //    pll_locked.export
		input  wire        sdcard_MISO,                //        sdcard.MISO
		output wire        sdcard_MOSI,                //              .MOSI
		output wire        sdcard_SCLK,                //              .SCLK
		output wire        sdcard_SS_n,                //              .SS_n
		input  wire [11:0] sw_export                   //            sw.export
	);

	wire         altpll_0_c0_clk;                                                                                     // altpll_0:c0 -> [addr_router:clk, addr_router_001:clk, addr_router_002:clk, addr_router_003:clk, burst_adapter:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_demux_002:clk, cmd_xbar_demux_003:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cmd_xbar_mux_002:clk, cmd_xbar_mux_013:clk, crosser:in_clk, crosser_001:out_clk, data_format_adapter:clk, fifo_0:wrclock, fifo_0_in_csr_translator:clk, fifo_0_in_csr_translator_avalon_universal_slave_0_agent:clk, fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, fifo_0_in_translator:clk, fifo_0_in_translator_avalon_universal_slave_0_agent:clk, fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, flash_0:clk, hexdisp_0:clk, hexdisp_0_ctrl_translator:clk, hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:clk, hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_005:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, id_router_009:clk, id_router_010:clk, id_router_011:clk, id_router_012:clk, id_router_013:clk, irq_mapper:clk, m2vdd_hx8347a_0:clk, m2vdd_hx8347a_0_ctrl_translator:clk, m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:clk, m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, m2vdd_hx8347a_0_fbuf_translator:clk, m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:clk, m2vdec_0:csi_clk, m2vdec_0_control_translator:clk, m2vdec_0_control_translator_avalon_universal_slave_0_agent:clk, m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, m2vdec_0_fbuf_translator:clk, m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:clk, nios2_qsys_0:clk, nios2_qsys_0_data_master_translator:clk, nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_0_instruction_master_translator:clk, nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_0_jtag_debug_module_translator:clk, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_0:clk, pio_0_s1_translator:clk, pio_0_s1_translator_avalon_universal_slave_0_agent:clk, pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, ram_0:clk, ram_0_s1_translator:clk, ram_0_s1_translator_avalon_universal_slave_0_agent:clk, ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rom_0:clk_clk, rom_0_uas_translator:clk, rom_0_uas_translator_avalon_universal_slave_0_agent:clk, rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_demux_009:clk, rsp_xbar_demux_010:clk, rsp_xbar_demux_011:clk, rsp_xbar_demux_012:clk, rsp_xbar_demux_013:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rst_controller_001:clk, sdram_0:clk, sdram_0_s1_translator:clk, sdram_0_s1_translator_avalon_universal_slave_0_agent:clk, sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, spi_0:clk, spi_0_spi_control_port_translator:clk, spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:clk, spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sysid_qsys_0:clock, sysid_qsys_0_control_slave_translator:clk, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:clk, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timer_0:clk, timer_0_s1_translator:clk, timer_0_s1_translator_avalon_universal_slave_0_agent:clk, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timing_adapter:clk, width_adapter:clk, width_adapter_001:clk]
	wire         rom_0_tcm_chipselect_n_out;                                                                          // rom_0:tcm_chipselect_n_out -> flash_0:tcs_tcm_chipselect_n_out
	wire         rom_0_tcm_grant;                                                                                     // flash_0:grant -> rom_0:tcm_grant
	wire         rom_0_tcm_data_outen;                                                                                // rom_0:tcm_data_outen -> flash_0:tcs_tcm_data_outen
	wire         rom_0_tcm_request;                                                                                   // rom_0:tcm_request -> flash_0:request
	wire  [15:0] rom_0_tcm_data_out;                                                                                  // rom_0:tcm_data_out -> flash_0:tcs_tcm_data_out
	wire         rom_0_tcm_write_n_out;                                                                               // rom_0:tcm_write_n_out -> flash_0:tcs_tcm_write_n_out
	wire  [21:0] rom_0_tcm_address_out;                                                                               // rom_0:tcm_address_out -> flash_0:tcs_tcm_address_out
	wire  [15:0] rom_0_tcm_data_in;                                                                                   // flash_0:tcs_tcm_data_in -> rom_0:tcm_data_in
	wire         rom_0_tcm_read_n_out;                                                                                // rom_0:tcm_read_n_out -> flash_0:tcs_tcm_read_n_out
	wire         altpll_0_c2_clk;                                                                                     // altpll_0:c2 -> m2vdd_hx8347a_0:lcd_clk
	wire         m2vdec_0_fptr_updated;                                                                               // m2vdec_0:coe_fptr_updated -> m2vdd_hx8347a_0:fptr_updated
	wire  [10:0] m2vdd_hx8347a_0_fptr_address;                                                                        // m2vdd_hx8347a_0:fptr_address -> m2vdec_0:coe_fptr_address
	wire         m2vdec_0_fptr_number;                                                                                // m2vdec_0:coe_fptr_number -> m2vdd_hx8347a_0:fptr_number
	wire         data_format_adapter_out_valid;                                                                       // data_format_adapter:out_valid -> m2vdec_0:asi_stream_valid
	wire   [7:0] data_format_adapter_out_data;                                                                        // data_format_adapter:out_data -> m2vdec_0:asi_stream_data
	wire         data_format_adapter_out_ready;                                                                       // m2vdec_0:asi_stream_ready -> data_format_adapter:out_ready
	wire         fifo_0_out_valid;                                                                                    // fifo_0:avalonst_source_valid -> timing_adapter:in_valid
	wire  [31:0] fifo_0_out_data;                                                                                     // fifo_0:avalonst_source_data -> timing_adapter:in_data
	wire         fifo_0_out_ready;                                                                                    // timing_adapter:in_ready -> fifo_0:avalonst_source_ready
	wire         timing_adapter_out_valid;                                                                            // timing_adapter:out_valid -> data_format_adapter:in_valid
	wire  [31:0] timing_adapter_out_data;                                                                             // timing_adapter:out_data -> data_format_adapter:in_data
	wire         timing_adapter_out_ready;                                                                            // data_format_adapter:in_ready -> timing_adapter:out_ready
	wire         nios2_qsys_0_instruction_master_waitrequest;                                                         // nios2_qsys_0_instruction_master_translator:av_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [24:0] nios2_qsys_0_instruction_master_address;                                                             // nios2_qsys_0:i_address -> nios2_qsys_0_instruction_master_translator:av_address
	wire         nios2_qsys_0_instruction_master_read;                                                                // nios2_qsys_0:i_read -> nios2_qsys_0_instruction_master_translator:av_read
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                                                            // nios2_qsys_0_instruction_master_translator:av_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                                                                // nios2_qsys_0_data_master_translator:av_waitrequest -> nios2_qsys_0:d_waitrequest
	wire  [31:0] nios2_qsys_0_data_master_writedata;                                                                  // nios2_qsys_0:d_writedata -> nios2_qsys_0_data_master_translator:av_writedata
	wire  [24:0] nios2_qsys_0_data_master_address;                                                                    // nios2_qsys_0:d_address -> nios2_qsys_0_data_master_translator:av_address
	wire         nios2_qsys_0_data_master_write;                                                                      // nios2_qsys_0:d_write -> nios2_qsys_0_data_master_translator:av_write
	wire         nios2_qsys_0_data_master_read;                                                                       // nios2_qsys_0:d_read -> nios2_qsys_0_data_master_translator:av_read
	wire  [31:0] nios2_qsys_0_data_master_readdata;                                                                   // nios2_qsys_0_data_master_translator:av_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_debugaccess;                                                                // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> nios2_qsys_0_data_master_translator:av_debugaccess
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                                                                 // nios2_qsys_0:d_byteenable -> nios2_qsys_0_data_master_translator:av_byteenable
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                             // nios2_qsys_0_jtag_debug_module_translator:av_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire   [8:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address;                               // nios2_qsys_0_jtag_debug_module_translator:av_address -> nios2_qsys_0:jtag_debug_module_address
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                            // nios2_qsys_0_jtag_debug_module_translator:av_chipselect -> nios2_qsys_0:jtag_debug_module_select
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write;                                 // nios2_qsys_0_jtag_debug_module_translator:av_write -> nios2_qsys_0:jtag_debug_module_write
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                              // nios2_qsys_0:jtag_debug_module_readdata -> nios2_qsys_0_jtag_debug_module_translator:av_readdata
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                         // nios2_qsys_0_jtag_debug_module_translator:av_begintransfer -> nios2_qsys_0:jtag_debug_module_begintransfer
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                           // nios2_qsys_0_jtag_debug_module_translator:av_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [3:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                            // nios2_qsys_0_jtag_debug_module_translator:av_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire  [31:0] ram_0_s1_translator_avalon_anti_slave_0_writedata;                                                   // ram_0_s1_translator:av_writedata -> ram_0:writedata
	wire  [10:0] ram_0_s1_translator_avalon_anti_slave_0_address;                                                     // ram_0_s1_translator:av_address -> ram_0:address
	wire         ram_0_s1_translator_avalon_anti_slave_0_chipselect;                                                  // ram_0_s1_translator:av_chipselect -> ram_0:chipselect
	wire         ram_0_s1_translator_avalon_anti_slave_0_clken;                                                       // ram_0_s1_translator:av_clken -> ram_0:clken
	wire         ram_0_s1_translator_avalon_anti_slave_0_write;                                                       // ram_0_s1_translator:av_write -> ram_0:write
	wire  [31:0] ram_0_s1_translator_avalon_anti_slave_0_readdata;                                                    // ram_0:readdata -> ram_0_s1_translator:av_readdata
	wire   [3:0] ram_0_s1_translator_avalon_anti_slave_0_byteenable;                                                  // ram_0_s1_translator:av_byteenable -> ram_0:byteenable
	wire         rom_0_uas_translator_avalon_anti_slave_0_waitrequest;                                                // rom_0:uas_waitrequest -> rom_0_uas_translator:av_waitrequest
	wire   [1:0] rom_0_uas_translator_avalon_anti_slave_0_burstcount;                                                 // rom_0_uas_translator:av_burstcount -> rom_0:uas_burstcount
	wire  [15:0] rom_0_uas_translator_avalon_anti_slave_0_writedata;                                                  // rom_0_uas_translator:av_writedata -> rom_0:uas_writedata
	wire  [21:0] rom_0_uas_translator_avalon_anti_slave_0_address;                                                    // rom_0_uas_translator:av_address -> rom_0:uas_address
	wire         rom_0_uas_translator_avalon_anti_slave_0_lock;                                                       // rom_0_uas_translator:av_lock -> rom_0:uas_lock
	wire         rom_0_uas_translator_avalon_anti_slave_0_write;                                                      // rom_0_uas_translator:av_write -> rom_0:uas_write
	wire         rom_0_uas_translator_avalon_anti_slave_0_read;                                                       // rom_0_uas_translator:av_read -> rom_0:uas_read
	wire  [15:0] rom_0_uas_translator_avalon_anti_slave_0_readdata;                                                   // rom_0:uas_readdata -> rom_0_uas_translator:av_readdata
	wire         rom_0_uas_translator_avalon_anti_slave_0_debugaccess;                                                // rom_0_uas_translator:av_debugaccess -> rom_0:uas_debugaccess
	wire         rom_0_uas_translator_avalon_anti_slave_0_readdatavalid;                                              // rom_0:uas_readdatavalid -> rom_0_uas_translator:av_readdatavalid
	wire   [1:0] rom_0_uas_translator_avalon_anti_slave_0_byteenable;                                                 // rom_0_uas_translator:av_byteenable -> rom_0:uas_byteenable
	wire         sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address;                                   // sysid_qsys_0_control_slave_translator:av_address -> sysid_qsys_0:address
	wire  [31:0] sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata;                                  // sysid_qsys_0:readdata -> sysid_qsys_0_control_slave_translator:av_readdata
	wire  [31:0] altpll_0_pll_slave_translator_avalon_anti_slave_0_writedata;                                         // altpll_0_pll_slave_translator:av_writedata -> altpll_0:writedata
	wire   [1:0] altpll_0_pll_slave_translator_avalon_anti_slave_0_address;                                           // altpll_0_pll_slave_translator:av_address -> altpll_0:address
	wire         altpll_0_pll_slave_translator_avalon_anti_slave_0_write;                                             // altpll_0_pll_slave_translator:av_write -> altpll_0:write
	wire         altpll_0_pll_slave_translator_avalon_anti_slave_0_read;                                              // altpll_0_pll_slave_translator:av_read -> altpll_0:read
	wire  [31:0] altpll_0_pll_slave_translator_avalon_anti_slave_0_readdata;                                          // altpll_0:readdata -> altpll_0_pll_slave_translator:av_readdata
	wire         fifo_0_in_translator_avalon_anti_slave_0_waitrequest;                                                // fifo_0:avalonmm_write_slave_waitrequest -> fifo_0_in_translator:av_waitrequest
	wire  [31:0] fifo_0_in_translator_avalon_anti_slave_0_writedata;                                                  // fifo_0_in_translator:av_writedata -> fifo_0:avalonmm_write_slave_writedata
	wire         fifo_0_in_translator_avalon_anti_slave_0_address;                                                    // fifo_0_in_translator:av_address -> fifo_0:avalonmm_write_slave_address
	wire         fifo_0_in_translator_avalon_anti_slave_0_write;                                                      // fifo_0_in_translator:av_write -> fifo_0:avalonmm_write_slave_write
	wire  [31:0] fifo_0_in_csr_translator_avalon_anti_slave_0_writedata;                                              // fifo_0_in_csr_translator:av_writedata -> fifo_0:wrclk_control_slave_writedata
	wire   [2:0] fifo_0_in_csr_translator_avalon_anti_slave_0_address;                                                // fifo_0_in_csr_translator:av_address -> fifo_0:wrclk_control_slave_address
	wire         fifo_0_in_csr_translator_avalon_anti_slave_0_write;                                                  // fifo_0_in_csr_translator:av_write -> fifo_0:wrclk_control_slave_write
	wire         fifo_0_in_csr_translator_avalon_anti_slave_0_read;                                                   // fifo_0_in_csr_translator:av_read -> fifo_0:wrclk_control_slave_read
	wire  [31:0] fifo_0_in_csr_translator_avalon_anti_slave_0_readdata;                                               // fifo_0:wrclk_control_slave_readdata -> fifo_0_in_csr_translator:av_readdata
	wire  [31:0] m2vdec_0_control_translator_avalon_anti_slave_0_writedata;                                           // m2vdec_0_control_translator:av_writedata -> m2vdec_0:avs_control_writedata
	wire         m2vdec_0_control_translator_avalon_anti_slave_0_address;                                             // m2vdec_0_control_translator:av_address -> m2vdec_0:avs_control_address
	wire         m2vdec_0_control_translator_avalon_anti_slave_0_write;                                               // m2vdec_0_control_translator:av_write -> m2vdec_0:avs_control_write
	wire         m2vdec_0_control_translator_avalon_anti_slave_0_read;                                                // m2vdec_0_control_translator:av_read -> m2vdec_0:avs_control_read
	wire  [31:0] m2vdec_0_control_translator_avalon_anti_slave_0_readdata;                                            // m2vdec_0:avs_control_readdata -> m2vdec_0_control_translator:av_readdata
	wire         m2vdec_0_control_translator_avalon_anti_slave_0_readdatavalid;                                       // m2vdec_0:avs_control_readdatavalid -> m2vdec_0_control_translator:av_readdatavalid
	wire  [31:0] hexdisp_0_ctrl_translator_avalon_anti_slave_0_writedata;                                             // hexdisp_0_ctrl_translator:av_writedata -> hexdisp_0:ctrl_writedata
	wire   [1:0] hexdisp_0_ctrl_translator_avalon_anti_slave_0_address;                                               // hexdisp_0_ctrl_translator:av_address -> hexdisp_0:ctrl_address
	wire         hexdisp_0_ctrl_translator_avalon_anti_slave_0_write;                                                 // hexdisp_0_ctrl_translator:av_write -> hexdisp_0:ctrl_write
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_anti_slave_0_waitrequest;                                     // m2vdd_hx8347a_0:ctrl_waitrequest -> m2vdd_hx8347a_0_ctrl_translator:av_waitrequest
	wire  [31:0] m2vdd_hx8347a_0_ctrl_translator_avalon_anti_slave_0_writedata;                                       // m2vdd_hx8347a_0_ctrl_translator:av_writedata -> m2vdd_hx8347a_0:ctrl_writedata
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_anti_slave_0_write;                                           // m2vdd_hx8347a_0_ctrl_translator:av_write -> m2vdd_hx8347a_0:ctrl_write
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_anti_slave_0_read;                                            // m2vdd_hx8347a_0_ctrl_translator:av_read -> m2vdd_hx8347a_0:ctrl_read
	wire  [31:0] m2vdd_hx8347a_0_ctrl_translator_avalon_anti_slave_0_readdata;                                        // m2vdd_hx8347a_0:ctrl_readdata -> m2vdd_hx8347a_0_ctrl_translator:av_readdata
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_anti_slave_0_readdatavalid;                                   // m2vdd_hx8347a_0:ctrl_readdatavalid -> m2vdd_hx8347a_0_ctrl_translator:av_readdatavalid
	wire  [15:0] timer_0_s1_translator_avalon_anti_slave_0_writedata;                                                 // timer_0_s1_translator:av_writedata -> timer_0:writedata
	wire   [2:0] timer_0_s1_translator_avalon_anti_slave_0_address;                                                   // timer_0_s1_translator:av_address -> timer_0:address
	wire         timer_0_s1_translator_avalon_anti_slave_0_chipselect;                                                // timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	wire         timer_0_s1_translator_avalon_anti_slave_0_write;                                                     // timer_0_s1_translator:av_write -> timer_0:write_n
	wire  [15:0] timer_0_s1_translator_avalon_anti_slave_0_readdata;                                                  // timer_0:readdata -> timer_0_s1_translator:av_readdata
	wire  [15:0] spi_0_spi_control_port_translator_avalon_anti_slave_0_writedata;                                     // spi_0_spi_control_port_translator:av_writedata -> spi_0:data_from_cpu
	wire   [2:0] spi_0_spi_control_port_translator_avalon_anti_slave_0_address;                                       // spi_0_spi_control_port_translator:av_address -> spi_0:mem_addr
	wire         spi_0_spi_control_port_translator_avalon_anti_slave_0_chipselect;                                    // spi_0_spi_control_port_translator:av_chipselect -> spi_0:spi_select
	wire         spi_0_spi_control_port_translator_avalon_anti_slave_0_write;                                         // spi_0_spi_control_port_translator:av_write -> spi_0:write_n
	wire         spi_0_spi_control_port_translator_avalon_anti_slave_0_read;                                          // spi_0_spi_control_port_translator:av_read -> spi_0:read_n
	wire  [15:0] spi_0_spi_control_port_translator_avalon_anti_slave_0_readdata;                                      // spi_0:data_to_cpu -> spi_0_spi_control_port_translator:av_readdata
	wire   [1:0] pio_0_s1_translator_avalon_anti_slave_0_address;                                                     // pio_0_s1_translator:av_address -> pio_0:address
	wire  [31:0] pio_0_s1_translator_avalon_anti_slave_0_readdata;                                                    // pio_0:readdata -> pio_0_s1_translator:av_readdata
	wire         m2vdd_hx8347a_0_fbuf_waitrequest;                                                                    // m2vdd_hx8347a_0_fbuf_translator:av_waitrequest -> m2vdd_hx8347a_0:fbuf_waitrequest
	wire  [15:0] m2vdd_hx8347a_0_fbuf_writedata;                                                                      // m2vdd_hx8347a_0:fbuf_writedata -> m2vdd_hx8347a_0_fbuf_translator:av_writedata
	wire  [22:0] m2vdd_hx8347a_0_fbuf_address;                                                                        // m2vdd_hx8347a_0:fbuf_address -> m2vdd_hx8347a_0_fbuf_translator:av_address
	wire         m2vdd_hx8347a_0_fbuf_write;                                                                          // m2vdd_hx8347a_0:fbuf_write -> m2vdd_hx8347a_0_fbuf_translator:av_write
	wire         m2vdd_hx8347a_0_fbuf_read;                                                                           // m2vdd_hx8347a_0:fbuf_read -> m2vdd_hx8347a_0_fbuf_translator:av_read
	wire  [15:0] m2vdd_hx8347a_0_fbuf_readdata;                                                                       // m2vdd_hx8347a_0_fbuf_translator:av_readdata -> m2vdd_hx8347a_0:fbuf_readdata
	wire         m2vdd_hx8347a_0_fbuf_readdatavalid;                                                                  // m2vdd_hx8347a_0_fbuf_translator:av_readdatavalid -> m2vdd_hx8347a_0:fbuf_readdatavalid
	wire         m2vdec_0_fbuf_waitrequest;                                                                           // m2vdec_0_fbuf_translator:av_waitrequest -> m2vdec_0:avm_fbuf_waitrequest
	wire  [15:0] m2vdec_0_fbuf_writedata;                                                                             // m2vdec_0:avm_fbuf_writedata -> m2vdec_0_fbuf_translator:av_writedata
	wire  [22:0] m2vdec_0_fbuf_address;                                                                               // m2vdec_0:avm_fbuf_address -> m2vdec_0_fbuf_translator:av_address
	wire         m2vdec_0_fbuf_write;                                                                                 // m2vdec_0:avm_fbuf_write -> m2vdec_0_fbuf_translator:av_write
	wire         m2vdec_0_fbuf_read;                                                                                  // m2vdec_0:avm_fbuf_read -> m2vdec_0_fbuf_translator:av_read
	wire  [15:0] m2vdec_0_fbuf_readdata;                                                                              // m2vdec_0_fbuf_translator:av_readdata -> m2vdec_0:avm_fbuf_readdata
	wire         m2vdec_0_fbuf_readdatavalid;                                                                         // m2vdec_0_fbuf_translator:av_readdatavalid -> m2vdec_0:avm_fbuf_readdatavalid
	wire         sdram_0_s1_translator_avalon_anti_slave_0_waitrequest;                                               // sdram_0:za_waitrequest -> sdram_0_s1_translator:av_waitrequest
	wire  [15:0] sdram_0_s1_translator_avalon_anti_slave_0_writedata;                                                 // sdram_0_s1_translator:av_writedata -> sdram_0:az_data
	wire  [21:0] sdram_0_s1_translator_avalon_anti_slave_0_address;                                                   // sdram_0_s1_translator:av_address -> sdram_0:az_addr
	wire         sdram_0_s1_translator_avalon_anti_slave_0_chipselect;                                                // sdram_0_s1_translator:av_chipselect -> sdram_0:az_cs
	wire         sdram_0_s1_translator_avalon_anti_slave_0_write;                                                     // sdram_0_s1_translator:av_write -> sdram_0:az_wr_n
	wire         sdram_0_s1_translator_avalon_anti_slave_0_read;                                                      // sdram_0_s1_translator:av_read -> sdram_0:az_rd_n
	wire  [15:0] sdram_0_s1_translator_avalon_anti_slave_0_readdata;                                                  // sdram_0:za_data -> sdram_0_s1_translator:av_readdata
	wire         sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid;                                             // sdram_0:za_valid -> sdram_0_s1_translator:av_readdatavalid
	wire   [1:0] sdram_0_s1_translator_avalon_anti_slave_0_byteenable;                                                // sdram_0_s1_translator:av_byteenable -> sdram_0:az_be_n
	wire         pio_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // pio_0_s1_translator:uav_waitrequest -> pio_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_0_s1_translator:uav_burstcount
	wire  [31:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_0_s1_translator:uav_writedata
	wire  [24:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_0_s1_translator:uav_address
	wire         pio_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_0_s1_translator:uav_write
	wire         pio_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_0_s1_translator:uav_lock
	wire         pio_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_0_s1_translator:uav_read
	wire  [31:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // pio_0_s1_translator:uav_readdata -> pio_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // pio_0_s1_translator:uav_readdatavalid -> pio_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         pio_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_0_s1_translator:uav_debugaccess
	wire   [3:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_0_s1_translator:uav_byteenable
	wire         pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [82:0] pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [82:0] pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         rom_0_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // rom_0_uas_translator:uav_waitrequest -> rom_0_uas_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [1:0] rom_0_uas_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // rom_0_uas_translator_avalon_universal_slave_0_agent:m0_burstcount -> rom_0_uas_translator:uav_burstcount
	wire  [15:0] rom_0_uas_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // rom_0_uas_translator_avalon_universal_slave_0_agent:m0_writedata -> rom_0_uas_translator:uav_writedata
	wire  [24:0] rom_0_uas_translator_avalon_universal_slave_0_agent_m0_address;                                      // rom_0_uas_translator_avalon_universal_slave_0_agent:m0_address -> rom_0_uas_translator:uav_address
	wire         rom_0_uas_translator_avalon_universal_slave_0_agent_m0_write;                                        // rom_0_uas_translator_avalon_universal_slave_0_agent:m0_write -> rom_0_uas_translator:uav_write
	wire         rom_0_uas_translator_avalon_universal_slave_0_agent_m0_lock;                                         // rom_0_uas_translator_avalon_universal_slave_0_agent:m0_lock -> rom_0_uas_translator:uav_lock
	wire         rom_0_uas_translator_avalon_universal_slave_0_agent_m0_read;                                         // rom_0_uas_translator_avalon_universal_slave_0_agent:m0_read -> rom_0_uas_translator:uav_read
	wire  [15:0] rom_0_uas_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // rom_0_uas_translator:uav_readdata -> rom_0_uas_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         rom_0_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // rom_0_uas_translator:uav_readdatavalid -> rom_0_uas_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         rom_0_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // rom_0_uas_translator_avalon_universal_slave_0_agent:m0_debugaccess -> rom_0_uas_translator:uav_debugaccess
	wire   [1:0] rom_0_uas_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // rom_0_uas_translator_avalon_universal_slave_0_agent:m0_byteenable -> rom_0_uas_translator:uav_byteenable
	wire         rom_0_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // rom_0_uas_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         rom_0_uas_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // rom_0_uas_translator_avalon_universal_slave_0_agent:rf_source_valid -> rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         rom_0_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // rom_0_uas_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [64:0] rom_0_uas_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // rom_0_uas_translator_avalon_universal_slave_0_agent:rf_source_data -> rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         rom_0_uas_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> rom_0_uas_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> rom_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> rom_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> rom_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [64:0] rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> rom_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // rom_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_ready -> rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         rom_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // rom_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> rom_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [15:0] rom_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // rom_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> rom_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         rom_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // rom_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> rom_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // spi_0_spi_control_port_translator:uav_waitrequest -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> spi_0_spi_control_port_translator:uav_burstcount
	wire  [31:0] spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata;                       // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> spi_0_spi_control_port_translator:uav_writedata
	wire  [24:0] spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address;                         // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_address -> spi_0_spi_control_port_translator:uav_address
	wire         spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write;                           // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_write -> spi_0_spi_control_port_translator:uav_write
	wire         spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock;                            // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> spi_0_spi_control_port_translator:uav_lock
	wire         spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read;                            // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_read -> spi_0_spi_control_port_translator:uav_read
	wire  [31:0] spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata;                        // spi_0_spi_control_port_translator:uav_readdata -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // spi_0_spi_control_port_translator:uav_readdatavalid -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> spi_0_spi_control_port_translator:uav_debugaccess
	wire   [3:0] spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> spi_0_spi_control_port_translator:uav_byteenable
	wire         spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [82:0] spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data;                     // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [82:0] spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // hexdisp_0_ctrl_translator:uav_waitrequest -> hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> hexdisp_0_ctrl_translator:uav_burstcount
	wire  [31:0] hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                               // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> hexdisp_0_ctrl_translator:uav_writedata
	wire  [24:0] hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                                 // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> hexdisp_0_ctrl_translator:uav_address
	wire         hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                                   // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> hexdisp_0_ctrl_translator:uav_write
	wire         hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                                    // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> hexdisp_0_ctrl_translator:uav_lock
	wire         hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                                    // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> hexdisp_0_ctrl_translator:uav_read
	wire  [31:0] hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                                // hexdisp_0_ctrl_translator:uav_readdata -> hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // hexdisp_0_ctrl_translator:uav_readdatavalid -> hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hexdisp_0_ctrl_translator:uav_debugaccess
	wire   [3:0] hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> hexdisp_0_ctrl_translator:uav_byteenable
	wire         hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [82:0] hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;                             // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [82:0] hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // m2vdec_0_control_translator:uav_waitrequest -> m2vdec_0_control_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // m2vdec_0_control_translator_avalon_universal_slave_0_agent:m0_burstcount -> m2vdec_0_control_translator:uav_burstcount
	wire  [31:0] m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_writedata;                             // m2vdec_0_control_translator_avalon_universal_slave_0_agent:m0_writedata -> m2vdec_0_control_translator:uav_writedata
	wire  [24:0] m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_address;                               // m2vdec_0_control_translator_avalon_universal_slave_0_agent:m0_address -> m2vdec_0_control_translator:uav_address
	wire         m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_write;                                 // m2vdec_0_control_translator_avalon_universal_slave_0_agent:m0_write -> m2vdec_0_control_translator:uav_write
	wire         m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_lock;                                  // m2vdec_0_control_translator_avalon_universal_slave_0_agent:m0_lock -> m2vdec_0_control_translator:uav_lock
	wire         m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_read;                                  // m2vdec_0_control_translator_avalon_universal_slave_0_agent:m0_read -> m2vdec_0_control_translator:uav_read
	wire  [31:0] m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_readdata;                              // m2vdec_0_control_translator:uav_readdata -> m2vdec_0_control_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // m2vdec_0_control_translator:uav_readdatavalid -> m2vdec_0_control_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // m2vdec_0_control_translator_avalon_universal_slave_0_agent:m0_debugaccess -> m2vdec_0_control_translator:uav_debugaccess
	wire   [3:0] m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // m2vdec_0_control_translator_avalon_universal_slave_0_agent:m0_byteenable -> m2vdec_0_control_translator:uav_byteenable
	wire         m2vdec_0_control_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // m2vdec_0_control_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         m2vdec_0_control_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // m2vdec_0_control_translator_avalon_universal_slave_0_agent:rf_source_valid -> m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         m2vdec_0_control_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // m2vdec_0_control_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [82:0] m2vdec_0_control_translator_avalon_universal_slave_0_agent_rf_source_data;                           // m2vdec_0_control_translator_avalon_universal_slave_0_agent:rf_source_data -> m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         m2vdec_0_control_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> m2vdec_0_control_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> m2vdec_0_control_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> m2vdec_0_control_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> m2vdec_0_control_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [82:0] m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> m2vdec_0_control_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // m2vdec_0_control_translator_avalon_universal_slave_0_agent:rf_sink_ready -> m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         m2vdec_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // m2vdec_0_control_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> m2vdec_0_control_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] m2vdec_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // m2vdec_0_control_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> m2vdec_0_control_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         m2vdec_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // m2vdec_0_control_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> m2vdec_0_control_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	wire  [24:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	wire   [3:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [82:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [82:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // ram_0_s1_translator:uav_waitrequest -> ram_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // ram_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ram_0_s1_translator:uav_burstcount
	wire  [31:0] ram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // ram_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ram_0_s1_translator:uav_writedata
	wire  [24:0] ram_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // ram_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> ram_0_s1_translator:uav_address
	wire         ram_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // ram_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> ram_0_s1_translator:uav_write
	wire         ram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // ram_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ram_0_s1_translator:uav_lock
	wire         ram_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // ram_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> ram_0_s1_translator:uav_read
	wire  [31:0] ram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // ram_0_s1_translator:uav_readdata -> ram_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // ram_0_s1_translator:uav_readdatavalid -> ram_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // ram_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ram_0_s1_translator:uav_debugaccess
	wire   [3:0] ram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // ram_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ram_0_s1_translator:uav_byteenable
	wire         ram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // ram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // ram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // ram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [82:0] ram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // ram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [82:0] ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // ram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // ram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] ram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // ram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // ram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // altpll_0_pll_slave_translator:uav_waitrequest -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> altpll_0_pll_slave_translator:uav_burstcount
	wire  [31:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                           // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> altpll_0_pll_slave_translator:uav_writedata
	wire  [24:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_address;                             // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_address -> altpll_0_pll_slave_translator:uav_address
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_write;                               // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_write -> altpll_0_pll_slave_translator:uav_write
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_lock -> altpll_0_pll_slave_translator:uav_lock
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_read;                                // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_read -> altpll_0_pll_slave_translator:uav_read
	wire  [31:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                            // altpll_0_pll_slave_translator:uav_readdata -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // altpll_0_pll_slave_translator:uav_readdatavalid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> altpll_0_pll_slave_translator:uav_debugaccess
	wire   [3:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> altpll_0_pll_slave_translator:uav_byteenable
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [82:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                         // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [82:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire  [31:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                   // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                    // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                   // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest;                           // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_data_master_translator:uav_waitrequest
	wire   [2:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount;                            // nios2_qsys_0_data_master_translator:uav_burstcount -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata;                             // nios2_qsys_0_data_master_translator:uav_writedata -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [24:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_address;                               // nios2_qsys_0_data_master_translator:uav_address -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock;                                  // nios2_qsys_0_data_master_translator:uav_lock -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_write;                                 // nios2_qsys_0_data_master_translator:uav_write -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_read;                                  // nios2_qsys_0_data_master_translator:uav_read -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata;                              // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_data_master_translator:uav_readdata
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess;                           // nios2_qsys_0_data_master_translator:uav_debugaccess -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable;                            // nios2_qsys_0_data_master_translator:uav_byteenable -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid;                         // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_data_master_translator:uav_readdatavalid
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // fifo_0_in_csr_translator:uav_waitrequest -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_0_in_csr_translator:uav_burstcount
	wire  [31:0] fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                                // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_0_in_csr_translator:uav_writedata
	wire  [24:0] fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                                  // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_0_in_csr_translator:uav_address
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                                    // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_0_in_csr_translator:uav_write
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                     // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_0_in_csr_translator:uav_lock
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                                     // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_0_in_csr_translator:uav_read
	wire  [31:0] fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // fifo_0_in_csr_translator:uav_readdata -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // fifo_0_in_csr_translator:uav_readdatavalid -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_0_in_csr_translator:uav_debugaccess
	wire   [3:0] fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_0_in_csr_translator:uav_byteenable
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [82:0] fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                              // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [82:0] fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest;                    // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_instruction_master_translator:uav_waitrequest
	wire   [2:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount;                     // nios2_qsys_0_instruction_master_translator:uav_burstcount -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata;                      // nios2_qsys_0_instruction_master_translator:uav_writedata -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [24:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address;                        // nios2_qsys_0_instruction_master_translator:uav_address -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock;                           // nios2_qsys_0_instruction_master_translator:uav_lock -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write;                          // nios2_qsys_0_instruction_master_translator:uav_write -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read;                           // nios2_qsys_0_instruction_master_translator:uav_read -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata;                       // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_instruction_master_translator:uav_readdata
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess;                    // nios2_qsys_0_instruction_master_translator:uav_debugaccess -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable;                     // nios2_qsys_0_instruction_master_translator:uav_byteenable -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid;                  // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_instruction_master_translator:uav_readdatavalid
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // sysid_qsys_0_control_slave_translator:uav_waitrequest -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_qsys_0_control_slave_translator:uav_burstcount
	wire  [31:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                   // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_qsys_0_control_slave_translator:uav_writedata
	wire  [24:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                     // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_qsys_0_control_slave_translator:uav_address
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                       // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_qsys_0_control_slave_translator:uav_write
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                        // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_qsys_0_control_slave_translator:uav_lock
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                        // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_qsys_0_control_slave_translator:uav_read
	wire  [31:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                    // sysid_qsys_0_control_slave_translator:uav_readdata -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // sysid_qsys_0_control_slave_translator:uav_readdatavalid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_qsys_0_control_slave_translator:uav_debugaccess
	wire   [3:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_qsys_0_control_slave_translator:uav_byteenable
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [82:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                 // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [82:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // m2vdd_hx8347a_0_ctrl_translator:uav_waitrequest -> m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> m2vdd_hx8347a_0_ctrl_translator:uav_burstcount
	wire  [31:0] m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                         // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> m2vdd_hx8347a_0_ctrl_translator:uav_writedata
	wire  [24:0] m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                           // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> m2vdd_hx8347a_0_ctrl_translator:uav_address
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                             // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> m2vdd_hx8347a_0_ctrl_translator:uav_write
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                              // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> m2vdd_hx8347a_0_ctrl_translator:uav_lock
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                              // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> m2vdd_hx8347a_0_ctrl_translator:uav_read
	wire  [31:0] m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                          // m2vdd_hx8347a_0_ctrl_translator:uav_readdata -> m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // m2vdd_hx8347a_0_ctrl_translator:uav_readdatavalid -> m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> m2vdd_hx8347a_0_ctrl_translator:uav_debugaccess
	wire   [3:0] m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> m2vdd_hx8347a_0_ctrl_translator:uav_byteenable
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [82:0] m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;                       // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [82:0] m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // nios2_qsys_0_jtag_debug_module_translator:uav_waitrequest -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_qsys_0_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;               // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_qsys_0_jtag_debug_module_translator:uav_writedata
	wire  [24:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                 // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_qsys_0_jtag_debug_module_translator:uav_address
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                   // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_qsys_0_jtag_debug_module_translator:uav_write
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_qsys_0_jtag_debug_module_translator:uav_lock
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_qsys_0_jtag_debug_module_translator:uav_read
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                // nios2_qsys_0_jtag_debug_module_translator:uav_readdata -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // nios2_qsys_0_jtag_debug_module_translator:uav_readdatavalid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_qsys_0_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_qsys_0_jtag_debug_module_translator:uav_byteenable
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;            // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [82:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;             // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;            // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [82:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // fifo_0_in_translator:uav_waitrequest -> fifo_0_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fifo_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // fifo_0_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_0_in_translator:uav_burstcount
	wire  [31:0] fifo_0_in_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // fifo_0_in_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_0_in_translator:uav_writedata
	wire  [24:0] fifo_0_in_translator_avalon_universal_slave_0_agent_m0_address;                                      // fifo_0_in_translator_avalon_universal_slave_0_agent:m0_address -> fifo_0_in_translator:uav_address
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_m0_write;                                        // fifo_0_in_translator_avalon_universal_slave_0_agent:m0_write -> fifo_0_in_translator:uav_write
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_m0_lock;                                         // fifo_0_in_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_0_in_translator:uav_lock
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_m0_read;                                         // fifo_0_in_translator_avalon_universal_slave_0_agent:m0_read -> fifo_0_in_translator:uav_read
	wire  [31:0] fifo_0_in_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // fifo_0_in_translator:uav_readdata -> fifo_0_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // fifo_0_in_translator:uav_readdatavalid -> fifo_0_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // fifo_0_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_0_in_translator:uav_debugaccess
	wire   [3:0] fifo_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // fifo_0_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_0_in_translator:uav_byteenable
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // fifo_0_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // fifo_0_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // fifo_0_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [82:0] fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // fifo_0_in_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_0_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_0_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_0_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_0_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [82:0] fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_0_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // fifo_0_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // fifo_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] fifo_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // fifo_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // fifo_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_0_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_waitrequest;                               // m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:av_waitrequest -> m2vdd_hx8347a_0_fbuf_translator:uav_waitrequest
	wire   [1:0] m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_burstcount;                                // m2vdd_hx8347a_0_fbuf_translator:uav_burstcount -> m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [15:0] m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_writedata;                                 // m2vdd_hx8347a_0_fbuf_translator:uav_writedata -> m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:av_writedata
	wire  [22:0] m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_address;                                   // m2vdd_hx8347a_0_fbuf_translator:uav_address -> m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:av_address
	wire         m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_lock;                                      // m2vdd_hx8347a_0_fbuf_translator:uav_lock -> m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:av_lock
	wire         m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_write;                                     // m2vdd_hx8347a_0_fbuf_translator:uav_write -> m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:av_write
	wire         m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_read;                                      // m2vdd_hx8347a_0_fbuf_translator:uav_read -> m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:av_read
	wire  [15:0] m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_readdata;                                  // m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:av_readdata -> m2vdd_hx8347a_0_fbuf_translator:uav_readdata
	wire         m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_debugaccess;                               // m2vdd_hx8347a_0_fbuf_translator:uav_debugaccess -> m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [1:0] m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_byteenable;                                // m2vdd_hx8347a_0_fbuf_translator:uav_byteenable -> m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:av_byteenable
	wire         m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_readdatavalid;                             // m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:av_readdatavalid -> m2vdd_hx8347a_0_fbuf_translator:uav_readdatavalid
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // sdram_0_s1_translator:uav_waitrequest -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [1:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_0_s1_translator:uav_burstcount
	wire  [15:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_0_s1_translator:uav_writedata
	wire  [22:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_0_s1_translator:uav_address
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_0_s1_translator:uav_write
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_0_s1_translator:uav_lock
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_0_s1_translator:uav_read
	wire  [15:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // sdram_0_s1_translator:uav_readdata -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // sdram_0_s1_translator:uav_readdatavalid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_0_s1_translator:uav_debugaccess
	wire   [1:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_0_s1_translator:uav_byteenable
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [54:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [54:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [15:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         m2vdec_0_fbuf_translator_avalon_universal_master_0_waitrequest;                                      // m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:av_waitrequest -> m2vdec_0_fbuf_translator:uav_waitrequest
	wire   [1:0] m2vdec_0_fbuf_translator_avalon_universal_master_0_burstcount;                                       // m2vdec_0_fbuf_translator:uav_burstcount -> m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [15:0] m2vdec_0_fbuf_translator_avalon_universal_master_0_writedata;                                        // m2vdec_0_fbuf_translator:uav_writedata -> m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:av_writedata
	wire  [22:0] m2vdec_0_fbuf_translator_avalon_universal_master_0_address;                                          // m2vdec_0_fbuf_translator:uav_address -> m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:av_address
	wire         m2vdec_0_fbuf_translator_avalon_universal_master_0_lock;                                             // m2vdec_0_fbuf_translator:uav_lock -> m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:av_lock
	wire         m2vdec_0_fbuf_translator_avalon_universal_master_0_write;                                            // m2vdec_0_fbuf_translator:uav_write -> m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:av_write
	wire         m2vdec_0_fbuf_translator_avalon_universal_master_0_read;                                             // m2vdec_0_fbuf_translator:uav_read -> m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:av_read
	wire  [15:0] m2vdec_0_fbuf_translator_avalon_universal_master_0_readdata;                                         // m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:av_readdata -> m2vdec_0_fbuf_translator:uav_readdata
	wire         m2vdec_0_fbuf_translator_avalon_universal_master_0_debugaccess;                                      // m2vdec_0_fbuf_translator:uav_debugaccess -> m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [1:0] m2vdec_0_fbuf_translator_avalon_universal_master_0_byteenable;                                       // m2vdec_0_fbuf_translator:uav_byteenable -> m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:av_byteenable
	wire         m2vdec_0_fbuf_translator_avalon_universal_master_0_readdatavalid;                                    // m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:av_readdatavalid -> m2vdec_0_fbuf_translator:uav_readdatavalid
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;           // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                 // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;         // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [81:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                  // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                 // addr_router:sink_ready -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                  // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid;                        // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [81:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data;                         // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready;                        // addr_router_001:sink_ready -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                   // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [81:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router:sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // ram_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         ram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // ram_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         ram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // ram_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [81:0] ram_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // ram_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         ram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_001:sink_ready -> ram_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         rom_0_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // rom_0_uas_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         rom_0_uas_translator_avalon_universal_slave_0_agent_rp_valid;                                        // rom_0_uas_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         rom_0_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // rom_0_uas_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [63:0] rom_0_uas_translator_avalon_universal_slave_0_agent_rp_data;                                         // rom_0_uas_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         rom_0_uas_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_002:sink_ready -> rom_0_uas_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                       // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [81:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                        // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router_003:sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid;                               // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [81:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_data;                                // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_004:sink_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // fifo_0_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rp_valid;                                        // fifo_0_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // fifo_0_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [81:0] fifo_0_in_translator_avalon_universal_slave_0_agent_rp_data;                                         // fifo_0_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         fifo_0_in_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_005:sink_ready -> fifo_0_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                    // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [81:0] fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                                     // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_006:sink_ready -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         m2vdec_0_control_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // m2vdec_0_control_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire         m2vdec_0_control_translator_avalon_universal_slave_0_agent_rp_valid;                                 // m2vdec_0_control_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire         m2vdec_0_control_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // m2vdec_0_control_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [81:0] m2vdec_0_control_translator_avalon_universal_slave_0_agent_rp_data;                                  // m2vdec_0_control_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire         m2vdec_0_control_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_007:sink_ready -> m2vdec_0_control_translator_avalon_universal_slave_0_agent:rp_ready
	wire         hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire         hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                                   // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire         hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [81:0] hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                                    // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire         hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_008:sink_ready -> hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                             // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [81:0] m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                              // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire         m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_009:sink_ready -> m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [81:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_010:sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire         spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid;                           // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire         spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [81:0] spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data;                            // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire         spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_011:sink_ready -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	wire         pio_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // pio_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire         pio_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // pio_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire         pio_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // pio_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [81:0] pio_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // pio_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire         pio_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_012:sink_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent_cp_endofpacket;                      // m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire         m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent_cp_valid;                            // m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire         m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent_cp_startofpacket;                    // m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [53:0] m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent_cp_data;                             // m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire         m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent_cp_ready;                            // addr_router_002:sink_ready -> m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:cp_ready
	wire         m2vdec_0_fbuf_translator_avalon_universal_master_0_agent_cp_endofpacket;                             // m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire         m2vdec_0_fbuf_translator_avalon_universal_master_0_agent_cp_valid;                                   // m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire         m2vdec_0_fbuf_translator_avalon_universal_master_0_agent_cp_startofpacket;                           // m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire  [53:0] m2vdec_0_fbuf_translator_avalon_universal_master_0_agent_cp_data;                                    // m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire         m2vdec_0_fbuf_translator_avalon_universal_master_0_agent_cp_ready;                                   // addr_router_003:sink_ready -> m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:cp_ready
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [53:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_013:sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         burst_adapter_source0_endofpacket;                                                                   // burst_adapter:source0_endofpacket -> rom_0_uas_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_source0_valid;                                                                         // burst_adapter:source0_valid -> rom_0_uas_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_source0_startofpacket;                                                                 // burst_adapter:source0_startofpacket -> rom_0_uas_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [63:0] burst_adapter_source0_data;                                                                          // burst_adapter:source0_data -> rom_0_uas_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_source0_ready;                                                                         // rom_0_uas_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire  [12:0] burst_adapter_source0_channel;                                                                       // burst_adapter:source0_channel -> rom_0_uas_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rst_controller_reset_out_reset;                                                                      // rst_controller:reset_out -> [altpll_0:reset, altpll_0_pll_slave_translator:reset, altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:reset, altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser:out_reset, crosser_001:in_reset, id_router_004:reset, rsp_xbar_demux_004:reset]
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                                                          // nios2_qsys_0:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in0]
	wire         rst_controller_001_reset_out_reset;                                                                  // rst_controller_001:reset_out -> [addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, burst_adapter:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_013:reset, crosser:in_reset, crosser_001:out_reset, data_format_adapter:reset_n, fifo_0:reset_n, fifo_0_in_csr_translator:reset, fifo_0_in_csr_translator_avalon_universal_slave_0_agent:reset, fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo_0_in_translator:reset, fifo_0_in_translator_avalon_universal_slave_0_agent:reset, fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, flash_0:reset, hexdisp_0:reset_n, hexdisp_0_ctrl_translator:reset, hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:reset, hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, irq_mapper:reset, m2vdd_hx8347a_0:reset_n, m2vdd_hx8347a_0_ctrl_translator:reset, m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:reset, m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, m2vdd_hx8347a_0_fbuf_translator:reset, m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:reset, m2vdec_0:rsi_reset_n, m2vdec_0_control_translator:reset, m2vdec_0_control_translator_avalon_universal_slave_0_agent:reset, m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, m2vdec_0_fbuf_translator:reset, m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0:reset_n, nios2_qsys_0_data_master_translator:reset, nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_instruction_master_translator:reset, nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_0:reset_n, pio_0_s1_translator:reset, pio_0_s1_translator_avalon_universal_slave_0_agent:reset, pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ram_0:reset, ram_0_s1_translator:reset, ram_0_s1_translator_avalon_universal_slave_0_agent:reset, ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rom_0:reset_reset, rom_0_uas_translator:reset, rom_0_uas_translator_avalon_universal_slave_0_agent:reset, rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, sdram_0:reset_n, sdram_0_s1_translator:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, spi_0:reset_n, spi_0_spi_control_port_translator:reset, spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:reset, spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid_qsys_0:reset_n, sysid_qsys_0_control_slave_translator:reset, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_0:reset_n, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timing_adapter:reset_n, width_adapter:reset, width_adapter_001:reset]
	wire         cmd_xbar_demux_src0_endofpacket;                                                                     // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                           // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                   // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [81:0] cmd_xbar_demux_src0_data;                                                                            // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire  [12:0] cmd_xbar_demux_src0_channel;                                                                         // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                           // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                     // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                           // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                   // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [81:0] cmd_xbar_demux_src1_data;                                                                            // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire  [12:0] cmd_xbar_demux_src1_channel;                                                                         // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                           // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_src2_endofpacket;                                                                     // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                                           // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                                   // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [81:0] cmd_xbar_demux_src2_data;                                                                            // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire  [12:0] cmd_xbar_demux_src2_channel;                                                                         // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire         cmd_xbar_demux_src2_ready;                                                                           // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                                 // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                       // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                               // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [81:0] cmd_xbar_demux_001_src0_data;                                                                        // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire  [12:0] cmd_xbar_demux_001_src0_channel;                                                                     // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                       // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                                 // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                       // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                               // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [81:0] cmd_xbar_demux_001_src1_data;                                                                        // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire  [12:0] cmd_xbar_demux_001_src1_channel;                                                                     // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                       // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                                 // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                       // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                               // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [81:0] cmd_xbar_demux_001_src2_data;                                                                        // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire  [12:0] cmd_xbar_demux_001_src2_channel;                                                                     // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire         cmd_xbar_demux_001_src2_ready;                                                                       // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                                 // cmd_xbar_demux_001:src3_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                                       // cmd_xbar_demux_001:src3_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                               // cmd_xbar_demux_001:src3_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [81:0] cmd_xbar_demux_001_src3_data;                                                                        // cmd_xbar_demux_001:src3_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] cmd_xbar_demux_001_src3_channel;                                                                     // cmd_xbar_demux_001:src3_channel -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src5_endofpacket;                                                                 // cmd_xbar_demux_001:src5_endofpacket -> fifo_0_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src5_valid;                                                                       // cmd_xbar_demux_001:src5_valid -> fifo_0_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src5_startofpacket;                                                               // cmd_xbar_demux_001:src5_startofpacket -> fifo_0_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [81:0] cmd_xbar_demux_001_src5_data;                                                                        // cmd_xbar_demux_001:src5_data -> fifo_0_in_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] cmd_xbar_demux_001_src5_channel;                                                                     // cmd_xbar_demux_001:src5_channel -> fifo_0_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src6_endofpacket;                                                                 // cmd_xbar_demux_001:src6_endofpacket -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src6_valid;                                                                       // cmd_xbar_demux_001:src6_valid -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src6_startofpacket;                                                               // cmd_xbar_demux_001:src6_startofpacket -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [81:0] cmd_xbar_demux_001_src6_data;                                                                        // cmd_xbar_demux_001:src6_data -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] cmd_xbar_demux_001_src6_channel;                                                                     // cmd_xbar_demux_001:src6_channel -> fifo_0_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src7_endofpacket;                                                                 // cmd_xbar_demux_001:src7_endofpacket -> m2vdec_0_control_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src7_valid;                                                                       // cmd_xbar_demux_001:src7_valid -> m2vdec_0_control_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src7_startofpacket;                                                               // cmd_xbar_demux_001:src7_startofpacket -> m2vdec_0_control_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [81:0] cmd_xbar_demux_001_src7_data;                                                                        // cmd_xbar_demux_001:src7_data -> m2vdec_0_control_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] cmd_xbar_demux_001_src7_channel;                                                                     // cmd_xbar_demux_001:src7_channel -> m2vdec_0_control_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src8_endofpacket;                                                                 // cmd_xbar_demux_001:src8_endofpacket -> hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src8_valid;                                                                       // cmd_xbar_demux_001:src8_valid -> hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src8_startofpacket;                                                               // cmd_xbar_demux_001:src8_startofpacket -> hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [81:0] cmd_xbar_demux_001_src8_data;                                                                        // cmd_xbar_demux_001:src8_data -> hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] cmd_xbar_demux_001_src8_channel;                                                                     // cmd_xbar_demux_001:src8_channel -> hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src9_endofpacket;                                                                 // cmd_xbar_demux_001:src9_endofpacket -> m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src9_valid;                                                                       // cmd_xbar_demux_001:src9_valid -> m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src9_startofpacket;                                                               // cmd_xbar_demux_001:src9_startofpacket -> m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [81:0] cmd_xbar_demux_001_src9_data;                                                                        // cmd_xbar_demux_001:src9_data -> m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] cmd_xbar_demux_001_src9_channel;                                                                     // cmd_xbar_demux_001:src9_channel -> m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src10_endofpacket;                                                                // cmd_xbar_demux_001:src10_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src10_valid;                                                                      // cmd_xbar_demux_001:src10_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src10_startofpacket;                                                              // cmd_xbar_demux_001:src10_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [81:0] cmd_xbar_demux_001_src10_data;                                                                       // cmd_xbar_demux_001:src10_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] cmd_xbar_demux_001_src10_channel;                                                                    // cmd_xbar_demux_001:src10_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src11_endofpacket;                                                                // cmd_xbar_demux_001:src11_endofpacket -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src11_valid;                                                                      // cmd_xbar_demux_001:src11_valid -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src11_startofpacket;                                                              // cmd_xbar_demux_001:src11_startofpacket -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [81:0] cmd_xbar_demux_001_src11_data;                                                                       // cmd_xbar_demux_001:src11_data -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] cmd_xbar_demux_001_src11_channel;                                                                    // cmd_xbar_demux_001:src11_channel -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src12_endofpacket;                                                                // cmd_xbar_demux_001:src12_endofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src12_valid;                                                                      // cmd_xbar_demux_001:src12_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src12_startofpacket;                                                              // cmd_xbar_demux_001:src12_startofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [81:0] cmd_xbar_demux_001_src12_data;                                                                       // cmd_xbar_demux_001:src12_data -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] cmd_xbar_demux_001_src12_channel;                                                                    // cmd_xbar_demux_001:src12_channel -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                                     // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                           // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                   // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [81:0] rsp_xbar_demux_src0_data;                                                                            // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire  [12:0] rsp_xbar_demux_src0_channel;                                                                         // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                           // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                     // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                           // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                   // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [81:0] rsp_xbar_demux_src1_data;                                                                            // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire  [12:0] rsp_xbar_demux_src1_channel;                                                                         // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                           // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                                 // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                       // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                               // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [81:0] rsp_xbar_demux_001_src0_data;                                                                        // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire  [12:0] rsp_xbar_demux_001_src0_channel;                                                                     // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                       // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                                 // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                       // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                               // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [81:0] rsp_xbar_demux_001_src1_data;                                                                        // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire  [12:0] rsp_xbar_demux_001_src1_channel;                                                                     // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                       // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                                 // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                       // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                               // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [81:0] rsp_xbar_demux_002_src0_data;                                                                        // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire  [12:0] rsp_xbar_demux_002_src0_channel;                                                                     // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                       // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_002_src1_endofpacket;                                                                 // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_002_src1_valid;                                                                       // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_002_src1_startofpacket;                                                               // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [81:0] rsp_xbar_demux_002_src1_data;                                                                        // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire  [12:0] rsp_xbar_demux_002_src1_channel;                                                                     // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_002_src1_ready;                                                                       // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                                 // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                       // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                               // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [81:0] rsp_xbar_demux_003_src0_data;                                                                        // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire  [12:0] rsp_xbar_demux_003_src0_channel;                                                                     // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                       // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                                 // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                       // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                               // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [81:0] rsp_xbar_demux_005_src0_data;                                                                        // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire  [12:0] rsp_xbar_demux_005_src0_channel;                                                                     // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                       // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                                 // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                                       // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                               // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [81:0] rsp_xbar_demux_006_src0_data;                                                                        // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire  [12:0] rsp_xbar_demux_006_src0_channel;                                                                     // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                                       // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         rsp_xbar_demux_007_src0_endofpacket;                                                                 // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire         rsp_xbar_demux_007_src0_valid;                                                                       // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire         rsp_xbar_demux_007_src0_startofpacket;                                                               // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [81:0] rsp_xbar_demux_007_src0_data;                                                                        // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire  [12:0] rsp_xbar_demux_007_src0_channel;                                                                     // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire         rsp_xbar_demux_007_src0_ready;                                                                       // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire         rsp_xbar_demux_008_src0_endofpacket;                                                                 // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire         rsp_xbar_demux_008_src0_valid;                                                                       // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire         rsp_xbar_demux_008_src0_startofpacket;                                                               // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [81:0] rsp_xbar_demux_008_src0_data;                                                                        // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire  [12:0] rsp_xbar_demux_008_src0_channel;                                                                     // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire         rsp_xbar_demux_008_src0_ready;                                                                       // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire         rsp_xbar_demux_009_src0_endofpacket;                                                                 // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire         rsp_xbar_demux_009_src0_valid;                                                                       // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire         rsp_xbar_demux_009_src0_startofpacket;                                                               // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [81:0] rsp_xbar_demux_009_src0_data;                                                                        // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire  [12:0] rsp_xbar_demux_009_src0_channel;                                                                     // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire         rsp_xbar_demux_009_src0_ready;                                                                       // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire         rsp_xbar_demux_010_src0_endofpacket;                                                                 // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire         rsp_xbar_demux_010_src0_valid;                                                                       // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	wire         rsp_xbar_demux_010_src0_startofpacket;                                                               // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [81:0] rsp_xbar_demux_010_src0_data;                                                                        // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	wire  [12:0] rsp_xbar_demux_010_src0_channel;                                                                     // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	wire         rsp_xbar_demux_010_src0_ready;                                                                       // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire         rsp_xbar_demux_011_src0_endofpacket;                                                                 // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire         rsp_xbar_demux_011_src0_valid;                                                                       // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	wire         rsp_xbar_demux_011_src0_startofpacket;                                                               // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [81:0] rsp_xbar_demux_011_src0_data;                                                                        // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	wire  [12:0] rsp_xbar_demux_011_src0_channel;                                                                     // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	wire         rsp_xbar_demux_011_src0_ready;                                                                       // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire         rsp_xbar_demux_012_src0_endofpacket;                                                                 // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire         rsp_xbar_demux_012_src0_valid;                                                                       // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink12_valid
	wire         rsp_xbar_demux_012_src0_startofpacket;                                                               // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [81:0] rsp_xbar_demux_012_src0_data;                                                                        // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink12_data
	wire  [12:0] rsp_xbar_demux_012_src0_channel;                                                                     // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink12_channel
	wire         rsp_xbar_demux_012_src0_ready;                                                                       // rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire         addr_router_src_endofpacket;                                                                         // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         addr_router_src_valid;                                                                               // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire         addr_router_src_startofpacket;                                                                       // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [81:0] addr_router_src_data;                                                                                // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire  [12:0] addr_router_src_channel;                                                                             // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire         addr_router_src_ready;                                                                               // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                        // rsp_xbar_mux:src_endofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                              // rsp_xbar_mux:src_valid -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                      // rsp_xbar_mux:src_startofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [81:0] rsp_xbar_mux_src_data;                                                                               // rsp_xbar_mux:src_data -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [12:0] rsp_xbar_mux_src_channel;                                                                            // rsp_xbar_mux:src_channel -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_src_ready;                                                                              // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire         addr_router_001_src_endofpacket;                                                                     // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         addr_router_001_src_valid;                                                                           // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire         addr_router_001_src_startofpacket;                                                                   // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [81:0] addr_router_001_src_data;                                                                            // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire  [12:0] addr_router_001_src_channel;                                                                         // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire         addr_router_001_src_ready;                                                                           // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                    // rsp_xbar_mux_001:src_endofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                          // rsp_xbar_mux_001:src_valid -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                                  // rsp_xbar_mux_001:src_startofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [81:0] rsp_xbar_mux_001_src_data;                                                                           // rsp_xbar_mux_001:src_data -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [12:0] rsp_xbar_mux_001_src_channel;                                                                        // rsp_xbar_mux_001:src_channel -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                          // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                        // cmd_xbar_mux:src_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                              // cmd_xbar_mux:src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                      // cmd_xbar_mux:src_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [81:0] cmd_xbar_mux_src_data;                                                                               // cmd_xbar_mux:src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] cmd_xbar_mux_src_channel;                                                                            // cmd_xbar_mux:src_channel -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                           // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                                 // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                         // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [81:0] id_router_src_data;                                                                                  // id_router:src_data -> rsp_xbar_demux:sink_data
	wire  [12:0] id_router_src_channel;                                                                               // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                                 // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                    // cmd_xbar_mux_001:src_endofpacket -> ram_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                          // cmd_xbar_mux_001:src_valid -> ram_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                                  // cmd_xbar_mux_001:src_startofpacket -> ram_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [81:0] cmd_xbar_mux_001_src_data;                                                                           // cmd_xbar_mux_001:src_data -> ram_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] cmd_xbar_mux_001_src_channel;                                                                        // cmd_xbar_mux_001:src_channel -> ram_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                          // ram_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire         id_router_001_src_endofpacket;                                                                       // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                             // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                                     // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [81:0] id_router_001_src_data;                                                                              // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire  [12:0] id_router_001_src_channel;                                                                           // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                             // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_demux_001_src3_ready;                                                                       // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire         id_router_003_src_endofpacket;                                                                       // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                             // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                     // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [81:0] id_router_003_src_data;                                                                              // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire  [12:0] id_router_003_src_channel;                                                                           // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                             // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         crosser_out_ready;                                                                                   // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser:out_ready
	wire         id_router_004_src_endofpacket;                                                                       // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                             // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                     // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [81:0] id_router_004_src_data;                                                                              // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire  [12:0] id_router_004_src_channel;                                                                           // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                             // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_demux_001_src5_ready;                                                                       // fifo_0_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire         id_router_005_src_endofpacket;                                                                       // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                             // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                     // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [81:0] id_router_005_src_data;                                                                              // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire  [12:0] id_router_005_src_channel;                                                                           // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                             // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_demux_001_src6_ready;                                                                       // fifo_0_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire         id_router_006_src_endofpacket;                                                                       // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         id_router_006_src_valid;                                                                             // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire         id_router_006_src_startofpacket;                                                                     // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [81:0] id_router_006_src_data;                                                                              // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire  [12:0] id_router_006_src_channel;                                                                           // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire         id_router_006_src_ready;                                                                             // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire         cmd_xbar_demux_001_src7_ready;                                                                       // m2vdec_0_control_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire         id_router_007_src_endofpacket;                                                                       // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire         id_router_007_src_valid;                                                                             // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire         id_router_007_src_startofpacket;                                                                     // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [81:0] id_router_007_src_data;                                                                              // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire  [12:0] id_router_007_src_channel;                                                                           // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire         id_router_007_src_ready;                                                                             // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire         cmd_xbar_demux_001_src8_ready;                                                                       // hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire         id_router_008_src_endofpacket;                                                                       // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire         id_router_008_src_valid;                                                                             // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire         id_router_008_src_startofpacket;                                                                     // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [81:0] id_router_008_src_data;                                                                              // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire  [12:0] id_router_008_src_channel;                                                                           // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire         id_router_008_src_ready;                                                                             // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire         cmd_xbar_demux_001_src9_ready;                                                                       // m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	wire         id_router_009_src_endofpacket;                                                                       // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire         id_router_009_src_valid;                                                                             // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire         id_router_009_src_startofpacket;                                                                     // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [81:0] id_router_009_src_data;                                                                              // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire  [12:0] id_router_009_src_channel;                                                                           // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire         id_router_009_src_ready;                                                                             // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire         cmd_xbar_demux_001_src10_ready;                                                                      // timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src10_ready
	wire         id_router_010_src_endofpacket;                                                                       // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire         id_router_010_src_valid;                                                                             // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire         id_router_010_src_startofpacket;                                                                     // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [81:0] id_router_010_src_data;                                                                              // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire  [12:0] id_router_010_src_channel;                                                                           // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire         id_router_010_src_ready;                                                                             // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire         cmd_xbar_demux_001_src11_ready;                                                                      // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src11_ready
	wire         id_router_011_src_endofpacket;                                                                       // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire         id_router_011_src_valid;                                                                             // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire         id_router_011_src_startofpacket;                                                                     // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [81:0] id_router_011_src_data;                                                                              // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire  [12:0] id_router_011_src_channel;                                                                           // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire         id_router_011_src_ready;                                                                             // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire         cmd_xbar_demux_001_src12_ready;                                                                      // pio_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src12_ready
	wire         id_router_012_src_endofpacket;                                                                       // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire         id_router_012_src_valid;                                                                             // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire         id_router_012_src_startofpacket;                                                                     // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [81:0] id_router_012_src_data;                                                                              // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire  [12:0] id_router_012_src_channel;                                                                           // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire         id_router_012_src_ready;                                                                             // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire         cmd_xbar_demux_002_src0_endofpacket;                                                                 // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_013:sink0_endofpacket
	wire         cmd_xbar_demux_002_src0_valid;                                                                       // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_013:sink0_valid
	wire         cmd_xbar_demux_002_src0_startofpacket;                                                               // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_013:sink0_startofpacket
	wire  [53:0] cmd_xbar_demux_002_src0_data;                                                                        // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_013:sink0_data
	wire   [1:0] cmd_xbar_demux_002_src0_channel;                                                                     // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_013:sink0_channel
	wire         cmd_xbar_demux_002_src0_ready;                                                                       // cmd_xbar_mux_013:sink0_ready -> cmd_xbar_demux_002:src0_ready
	wire         cmd_xbar_demux_003_src0_endofpacket;                                                                 // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_013:sink1_endofpacket
	wire         cmd_xbar_demux_003_src0_valid;                                                                       // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_013:sink1_valid
	wire         cmd_xbar_demux_003_src0_startofpacket;                                                               // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_013:sink1_startofpacket
	wire  [53:0] cmd_xbar_demux_003_src0_data;                                                                        // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_013:sink1_data
	wire   [1:0] cmd_xbar_demux_003_src0_channel;                                                                     // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_013:sink1_channel
	wire         cmd_xbar_demux_003_src0_ready;                                                                       // cmd_xbar_mux_013:sink1_ready -> cmd_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_013_src0_endofpacket;                                                                 // rsp_xbar_demux_013:src0_endofpacket -> m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_demux_013_src0_valid;                                                                       // rsp_xbar_demux_013:src0_valid -> m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_demux_013_src0_startofpacket;                                                               // rsp_xbar_demux_013:src0_startofpacket -> m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [53:0] rsp_xbar_demux_013_src0_data;                                                                        // rsp_xbar_demux_013:src0_data -> m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:rp_data
	wire   [1:0] rsp_xbar_demux_013_src0_channel;                                                                     // rsp_xbar_demux_013:src0_channel -> m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_demux_013_src1_endofpacket;                                                                 // rsp_xbar_demux_013:src1_endofpacket -> m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_demux_013_src1_valid;                                                                       // rsp_xbar_demux_013:src1_valid -> m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_demux_013_src1_startofpacket;                                                               // rsp_xbar_demux_013:src1_startofpacket -> m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [53:0] rsp_xbar_demux_013_src1_data;                                                                        // rsp_xbar_demux_013:src1_data -> m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:rp_data
	wire   [1:0] rsp_xbar_demux_013_src1_channel;                                                                     // rsp_xbar_demux_013:src1_channel -> m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:rp_channel
	wire         addr_router_002_src_endofpacket;                                                                     // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire         addr_router_002_src_valid;                                                                           // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire         addr_router_002_src_startofpacket;                                                                   // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [53:0] addr_router_002_src_data;                                                                            // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire   [1:0] addr_router_002_src_channel;                                                                         // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire         addr_router_002_src_ready;                                                                           // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire         rsp_xbar_demux_013_src0_ready;                                                                       // m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_013:src0_ready
	wire         addr_router_003_src_endofpacket;                                                                     // addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire         addr_router_003_src_valid;                                                                           // addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	wire         addr_router_003_src_startofpacket;                                                                   // addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire  [53:0] addr_router_003_src_data;                                                                            // addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	wire   [1:0] addr_router_003_src_channel;                                                                         // addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	wire         addr_router_003_src_ready;                                                                           // cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	wire         rsp_xbar_demux_013_src1_ready;                                                                       // m2vdec_0_fbuf_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_013:src1_ready
	wire         cmd_xbar_mux_013_src_endofpacket;                                                                    // cmd_xbar_mux_013:src_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_013_src_valid;                                                                          // cmd_xbar_mux_013:src_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_013_src_startofpacket;                                                                  // cmd_xbar_mux_013:src_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [53:0] cmd_xbar_mux_013_src_data;                                                                           // cmd_xbar_mux_013:src_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [1:0] cmd_xbar_mux_013_src_channel;                                                                        // cmd_xbar_mux_013:src_channel -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_013_src_ready;                                                                          // sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_013:src_ready
	wire         id_router_013_src_endofpacket;                                                                       // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire         id_router_013_src_valid;                                                                             // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire         id_router_013_src_startofpacket;                                                                     // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [53:0] id_router_013_src_data;                                                                              // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [1:0] id_router_013_src_channel;                                                                           // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire         id_router_013_src_ready;                                                                             // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire         cmd_xbar_mux_002_src_endofpacket;                                                                    // cmd_xbar_mux_002:src_endofpacket -> width_adapter:in_endofpacket
	wire         cmd_xbar_mux_002_src_valid;                                                                          // cmd_xbar_mux_002:src_valid -> width_adapter:in_valid
	wire         cmd_xbar_mux_002_src_startofpacket;                                                                  // cmd_xbar_mux_002:src_startofpacket -> width_adapter:in_startofpacket
	wire  [81:0] cmd_xbar_mux_002_src_data;                                                                           // cmd_xbar_mux_002:src_data -> width_adapter:in_data
	wire  [12:0] cmd_xbar_mux_002_src_channel;                                                                        // cmd_xbar_mux_002:src_channel -> width_adapter:in_channel
	wire         cmd_xbar_mux_002_src_ready;                                                                          // width_adapter:in_ready -> cmd_xbar_mux_002:src_ready
	wire         width_adapter_src_endofpacket;                                                                       // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire         width_adapter_src_valid;                                                                             // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire         width_adapter_src_startofpacket;                                                                     // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire  [63:0] width_adapter_src_data;                                                                              // width_adapter:out_data -> burst_adapter:sink0_data
	wire         width_adapter_src_ready;                                                                             // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire  [12:0] width_adapter_src_channel;                                                                           // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire         id_router_002_src_endofpacket;                                                                       // id_router_002:src_endofpacket -> width_adapter_001:in_endofpacket
	wire         id_router_002_src_valid;                                                                             // id_router_002:src_valid -> width_adapter_001:in_valid
	wire         id_router_002_src_startofpacket;                                                                     // id_router_002:src_startofpacket -> width_adapter_001:in_startofpacket
	wire  [63:0] id_router_002_src_data;                                                                              // id_router_002:src_data -> width_adapter_001:in_data
	wire  [12:0] id_router_002_src_channel;                                                                           // id_router_002:src_channel -> width_adapter_001:in_channel
	wire         id_router_002_src_ready;                                                                             // width_adapter_001:in_ready -> id_router_002:src_ready
	wire         width_adapter_001_src_endofpacket;                                                                   // width_adapter_001:out_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         width_adapter_001_src_valid;                                                                         // width_adapter_001:out_valid -> rsp_xbar_demux_002:sink_valid
	wire         width_adapter_001_src_startofpacket;                                                                 // width_adapter_001:out_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [81:0] width_adapter_001_src_data;                                                                          // width_adapter_001:out_data -> rsp_xbar_demux_002:sink_data
	wire         width_adapter_001_src_ready;                                                                         // rsp_xbar_demux_002:sink_ready -> width_adapter_001:out_ready
	wire  [12:0] width_adapter_001_src_channel;                                                                       // width_adapter_001:out_channel -> rsp_xbar_demux_002:sink_channel
	wire         crosser_out_endofpacket;                                                                             // crosser:out_endofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         crosser_out_valid;                                                                                   // crosser:out_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         crosser_out_startofpacket;                                                                           // crosser:out_startofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [81:0] crosser_out_data;                                                                                    // crosser:out_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] crosser_out_channel;                                                                                 // crosser:out_channel -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src4_endofpacket;                                                                 // cmd_xbar_demux_001:src4_endofpacket -> crosser:in_endofpacket
	wire         cmd_xbar_demux_001_src4_valid;                                                                       // cmd_xbar_demux_001:src4_valid -> crosser:in_valid
	wire         cmd_xbar_demux_001_src4_startofpacket;                                                               // cmd_xbar_demux_001:src4_startofpacket -> crosser:in_startofpacket
	wire  [81:0] cmd_xbar_demux_001_src4_data;                                                                        // cmd_xbar_demux_001:src4_data -> crosser:in_data
	wire  [12:0] cmd_xbar_demux_001_src4_channel;                                                                     // cmd_xbar_demux_001:src4_channel -> crosser:in_channel
	wire         cmd_xbar_demux_001_src4_ready;                                                                       // crosser:in_ready -> cmd_xbar_demux_001:src4_ready
	wire         crosser_001_out_endofpacket;                                                                         // crosser_001:out_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire         crosser_001_out_valid;                                                                               // crosser_001:out_valid -> rsp_xbar_mux_001:sink4_valid
	wire         crosser_001_out_startofpacket;                                                                       // crosser_001:out_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [81:0] crosser_001_out_data;                                                                                // crosser_001:out_data -> rsp_xbar_mux_001:sink4_data
	wire  [12:0] crosser_001_out_channel;                                                                             // crosser_001:out_channel -> rsp_xbar_mux_001:sink4_channel
	wire         crosser_001_out_ready;                                                                               // rsp_xbar_mux_001:sink4_ready -> crosser_001:out_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                                 // rsp_xbar_demux_004:src0_endofpacket -> crosser_001:in_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                       // rsp_xbar_demux_004:src0_valid -> crosser_001:in_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                               // rsp_xbar_demux_004:src0_startofpacket -> crosser_001:in_startofpacket
	wire  [81:0] rsp_xbar_demux_004_src0_data;                                                                        // rsp_xbar_demux_004:src0_data -> crosser_001:in_data
	wire  [12:0] rsp_xbar_demux_004_src0_channel;                                                                     // rsp_xbar_demux_004:src0_channel -> crosser_001:in_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                       // crosser_001:in_ready -> rsp_xbar_demux_004:src0_ready
	wire         irq_mapper_receiver0_irq;                                                                            // m2vdec_0:ins_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                                            // fifo_0:wrclk_control_slave_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                                            // timer_0:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                                            // spi_0:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                                                              // irq_mapper:sender_irq -> nios2_qsys_0:d_irq

	demo_de0_sys_altpll_0 altpll_0 (
		.clk       (clk_clk),                                                     //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),                              // inclk_interface_reset.reset
		.read      (altpll_0_pll_slave_translator_avalon_anti_slave_0_read),      //             pll_slave.read
		.write     (altpll_0_pll_slave_translator_avalon_anti_slave_0_write),     //                      .write
		.address   (altpll_0_pll_slave_translator_avalon_anti_slave_0_address),   //                      .address
		.readdata  (altpll_0_pll_slave_translator_avalon_anti_slave_0_readdata),  //                      .readdata
		.writedata (altpll_0_pll_slave_translator_avalon_anti_slave_0_writedata), //                      .writedata
		.c0        (altpll_0_c0_clk),                                             //                    c0.clk
		.c1        (sdrclk_clk),                                                  //                    c1.clk
		.c2        (altpll_0_c2_clk),                                             //                    c2.clk
		.areset    (pll_areset_export),                                           //        areset_conduit.export
		.locked    (pll_locked_export),                                           //        locked_conduit.export
		.phasedone (pll_phasedone_export)                                         //     phasedone_conduit.export
	);

	demo_de0_sys_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (altpll_0_c0_clk),                                                             //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                                         //                   reset_n.reset_n
		.d_address                             (nios2_qsys_0_data_master_address),                                            //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                               //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                                              //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                                        //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                                 //                          .waitrequest
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                             // custom_instruction_master.readra
	);

	demo_de0_sys_sysid_qsys_0 sysid_qsys_0 (
		.clock    (altpll_0_c0_clk),                                                    //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                                //         reset.reset_n
		.readdata (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	demo_de0_sys_ram_0 ram_0 (
		.clk        (altpll_0_c0_clk),                                    //   clk1.clk
		.address    (ram_0_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (ram_0_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (ram_0_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (ram_0_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (ram_0_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (ram_0_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (ram_0_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset)                  // reset1.reset
	);

	demo_de0_sys_rom_0 #(
		.TCM_ADDRESS_W                  (22),
		.TCM_DATA_W                     (16),
		.TCM_BYTEENABLE_W               (2),
		.TCM_READ_WAIT                  (70),
		.TCM_WRITE_WAIT                 (70),
		.TCM_SETUP_WAIT                 (35),
		.TCM_DATA_HOLD                  (0),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (2),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) rom_0 (
		.clk_clk              (altpll_0_c0_clk),                                        //   clk.clk
		.reset_reset          (rst_controller_001_reset_out_reset),                     // reset.reset
		.uas_address          (rom_0_uas_translator_avalon_anti_slave_0_address),       //   uas.address
		.uas_burstcount       (rom_0_uas_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.uas_read             (rom_0_uas_translator_avalon_anti_slave_0_read),          //      .read
		.uas_write            (rom_0_uas_translator_avalon_anti_slave_0_write),         //      .write
		.uas_waitrequest      (rom_0_uas_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (rom_0_uas_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.uas_byteenable       (rom_0_uas_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.uas_readdata         (rom_0_uas_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.uas_writedata        (rom_0_uas_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.uas_lock             (rom_0_uas_translator_avalon_anti_slave_0_lock),          //      .lock
		.uas_debugaccess      (rom_0_uas_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (rom_0_tcm_write_n_out),                                  //   tcm.write_n_out
		.tcm_read_n_out       (rom_0_tcm_read_n_out),                                   //      .read_n_out
		.tcm_chipselect_n_out (rom_0_tcm_chipselect_n_out),                             //      .chipselect_n_out
		.tcm_request          (rom_0_tcm_request),                                      //      .request
		.tcm_grant            (rom_0_tcm_grant),                                        //      .grant
		.tcm_address_out      (rom_0_tcm_address_out),                                  //      .address_out
		.tcm_data_out         (rom_0_tcm_data_out),                                     //      .data_out
		.tcm_data_outen       (rom_0_tcm_data_outen),                                   //      .data_outen
		.tcm_data_in          (rom_0_tcm_data_in)                                       //      .data_in
	);

	demo_de0_sys_flash_0 flash_0 (
		.clk                      (altpll_0_c0_clk),                    //   clk.clk
		.reset                    (rst_controller_001_reset_out_reset), // reset.reset
		.request                  (rom_0_tcm_request),                  //   tcs.request
		.grant                    (rom_0_tcm_grant),                    //      .grant
		.tcs_tcm_address_out      (rom_0_tcm_address_out),              //      .address_out
		.tcs_tcm_read_n_out       (rom_0_tcm_read_n_out),               //      .read_n_out
		.tcs_tcm_write_n_out      (rom_0_tcm_write_n_out),              //      .write_n_out
		.tcs_tcm_data_out         (rom_0_tcm_data_out),                 //      .data_out
		.tcs_tcm_data_outen       (rom_0_tcm_data_outen),               //      .data_outen
		.tcs_tcm_data_in          (rom_0_tcm_data_in),                  //      .data_in
		.tcs_tcm_chipselect_n_out (rom_0_tcm_chipselect_n_out),         //      .chipselect_n_out
		.tcm_address_out          (flash_tcm_address_out),              //   out.tcm_address_out
		.tcm_read_n_out           (flash_tcm_read_n_out),               //      .tcm_read_n_out
		.tcm_write_n_out          (flash_tcm_write_n_out),              //      .tcm_write_n_out
		.tcm_data_out             (flash_tcm_data_out),                 //      .tcm_data_out
		.tcm_chipselect_n_out     (flash_tcm_chipselect_n_out)          //      .tcm_chipselect_n_out
	);

	demo_de0_sys_fifo_0 fifo_0 (
		.wrclock                          (altpll_0_c0_clk),                                        //   clk_in.clk
		.reset_n                          (~rst_controller_001_reset_out_reset),                    // reset_in.reset_n
		.avalonmm_write_slave_writedata   (fifo_0_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (fifo_0_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_address     (fifo_0_in_translator_avalon_anti_slave_0_address),       //         .address
		.avalonmm_write_slave_waitrequest (fifo_0_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (fifo_0_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (fifo_0_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (fifo_0_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (fifo_0_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (fifo_0_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver1_irq),                               //   in_irq.irq
		.avalonst_source_valid            (fifo_0_out_valid),                                       //      out.valid
		.avalonst_source_data             (fifo_0_out_data),                                        //         .data
		.avalonst_source_ready            (fifo_0_out_ready)                                        //         .ready
	);

	m2vdec #(
		.MEM_WIDTH (23),
		.MVH_WIDTH (16),
		.MVV_WIDTH (15),
		.MBX_WIDTH (6),
		.MBY_WIDTH (5),
		.MBX_ADDER (6)
	) m2vdec_0 (
		.csi_clk                   (altpll_0_c0_clk),                                               //   clock.clk
		.rsi_reset_n               (~rst_controller_001_reset_out_reset),                           //   reset.reset_n
		.avs_control_address       (m2vdec_0_control_translator_avalon_anti_slave_0_address),       // control.address
		.avs_control_read          (m2vdec_0_control_translator_avalon_anti_slave_0_read),          //        .read
		.avs_control_readdata      (m2vdec_0_control_translator_avalon_anti_slave_0_readdata),      //        .readdata
		.avs_control_write         (m2vdec_0_control_translator_avalon_anti_slave_0_write),         //        .write
		.avs_control_writedata     (m2vdec_0_control_translator_avalon_anti_slave_0_writedata),     //        .writedata
		.avs_control_readdatavalid (m2vdec_0_control_translator_avalon_anti_slave_0_readdatavalid), //        .readdatavalid
		.ins_irq                   (irq_mapper_receiver0_irq),                                      //     irq.irq
		.asi_stream_data           (data_format_adapter_out_data),                                  //  stream.data
		.asi_stream_ready          (data_format_adapter_out_ready),                                 //        .ready
		.asi_stream_valid          (data_format_adapter_out_valid),                                 //        .valid
		.avm_fbuf_address          (m2vdec_0_fbuf_address),                                         //    fbuf.address
		.avm_fbuf_read             (m2vdec_0_fbuf_read),                                            //        .read
		.avm_fbuf_readdata         (m2vdec_0_fbuf_readdata),                                        //        .readdata
		.avm_fbuf_write            (m2vdec_0_fbuf_write),                                           //        .write
		.avm_fbuf_writedata        (m2vdec_0_fbuf_writedata),                                       //        .writedata
		.avm_fbuf_waitrequest      (m2vdec_0_fbuf_waitrequest),                                     //        .waitrequest
		.avm_fbuf_readdatavalid    (m2vdec_0_fbuf_readdatavalid),                                   //        .readdatavalid
		.coe_fptr_address          (m2vdd_hx8347a_0_fptr_address),                                  //    fptr.export
		.coe_fptr_updated          (m2vdec_0_fptr_updated),                                         //        .export
		.coe_fptr_number           (m2vdec_0_fptr_number)                                           //        .export
	);

	seg7led_static #(
		.DIGITS     (4),
		.ACTIVE_LOW (0)
	) hexdisp_0 (
		.clk            (altpll_0_c0_clk),                                         //  clock.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                     //  reset.reset_n
		.ctrl_address   (hexdisp_0_ctrl_translator_avalon_anti_slave_0_address),   //   ctrl.address
		.ctrl_write     (hexdisp_0_ctrl_translator_avalon_anti_slave_0_write),     //       .write
		.ctrl_writedata (hexdisp_0_ctrl_translator_avalon_anti_slave_0_writedata), //       .writedata
		.seg_a          (hd_a),                                                    // output.export
		.seg_b          (hd_b),                                                    //       .export
		.seg_c          (hd_c),                                                    //       .export
		.seg_d          (hd_d),                                                    //       .export
		.seg_e          (hd_e),                                                    //       .export
		.seg_f          (hd_f),                                                    //       .export
		.seg_g          (hd_g),                                                    //       .export
		.seg_dp         (hd_dp)                                                    //       .export
	);

	m2vdd_hx8347a #(
		.MEM_WIDTH (23),
		.MBX_WIDTH (6),
		.MBY_WIDTH (5)
	) m2vdd_hx8347a_0 (
		.clk                (altpll_0_c0_clk),                                                   //   clock.clk
		.reset_n            (~rst_controller_001_reset_out_reset),                               //   reset.reset_n
		.ctrl_read          (m2vdd_hx8347a_0_ctrl_translator_avalon_anti_slave_0_read),          //    ctrl.read
		.ctrl_readdata      (m2vdd_hx8347a_0_ctrl_translator_avalon_anti_slave_0_readdata),      //        .readdata
		.ctrl_write         (m2vdd_hx8347a_0_ctrl_translator_avalon_anti_slave_0_write),         //        .write
		.ctrl_writedata     (m2vdd_hx8347a_0_ctrl_translator_avalon_anti_slave_0_writedata),     //        .writedata
		.ctrl_waitrequest   (m2vdd_hx8347a_0_ctrl_translator_avalon_anti_slave_0_waitrequest),   //        .waitrequest
		.ctrl_readdatavalid (m2vdd_hx8347a_0_ctrl_translator_avalon_anti_slave_0_readdatavalid), //        .readdatavalid
		.lcd_clk            (altpll_0_c2_clk),                                                   // lcd_clk.clk
		.lcd_reset_n        (lcd_reset_n),                                                       //     lcd.export
		.lcd_cs             (lcd_cs),                                                            //        .export
		.lcd_rs             (lcd_rs),                                                            //        .export
		.lcd_data           (lcd_data),                                                          //        .export
		.lcd_write_n        (lcd_write_n),                                                       //        .export
		.lcd_read_n         (lcd_read_n),                                                        //        .export
		.fbuf_address       (m2vdd_hx8347a_0_fbuf_address),                                      //    fbuf.address
		.fbuf_read          (m2vdd_hx8347a_0_fbuf_read),                                         //        .read
		.fbuf_readdata      (m2vdd_hx8347a_0_fbuf_readdata),                                     //        .readdata
		.fbuf_write         (m2vdd_hx8347a_0_fbuf_write),                                        //        .write
		.fbuf_writedata     (m2vdd_hx8347a_0_fbuf_writedata),                                    //        .writedata
		.fbuf_waitrequest   (m2vdd_hx8347a_0_fbuf_waitrequest),                                  //        .waitrequest
		.fbuf_readdatavalid (m2vdd_hx8347a_0_fbuf_readdatavalid),                                //        .readdatavalid
		.fptr_address       (m2vdd_hx8347a_0_fptr_address),                                      //    fptr.export
		.fptr_updated       (m2vdec_0_fptr_updated),                                             //        .export
		.fptr_number        (m2vdec_0_fptr_number)                                               //        .export
	);

	demo_de0_sys_sdram_0 sdram_0 (
		.clk            (altpll_0_c0_clk),                                         //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                     // reset.reset_n
		.az_addr        (sdram_0_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_0_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_0_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_0_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_0_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_0_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_0_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_0_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdr_addr),                                                //  wire.export
		.zs_ba          (sdr_ba),                                                  //      .export
		.zs_cas_n       (sdr_cas_n),                                               //      .export
		.zs_cke         (sdr_cke),                                                 //      .export
		.zs_cs_n        (sdr_cs_n),                                                //      .export
		.zs_dq          (sdr_dq),                                                  //      .export
		.zs_dqm         (sdr_dqm),                                                 //      .export
		.zs_ras_n       (sdr_ras_n),                                               //      .export
		.zs_we_n        (sdr_we_n)                                                 //      .export
	);

	demo_de0_sys_data_format_adapter data_format_adapter (
		.clk       (altpll_0_c0_clk),                     //   clk.clk
		.reset_n   (~rst_controller_001_reset_out_reset), // reset.reset_n
		.in_ready  (timing_adapter_out_ready),            //    in.ready
		.in_valid  (timing_adapter_out_valid),            //      .valid
		.in_data   (timing_adapter_out_data),             //      .data
		.out_ready (data_format_adapter_out_ready),       //   out.ready
		.out_valid (data_format_adapter_out_valid),       //      .valid
		.out_data  (data_format_adapter_out_data)         //      .data
	);

	demo_de0_sys_timing_adapter timing_adapter (
		.clk       (altpll_0_c0_clk),                     //   clk.clk
		.reset_n   (~rst_controller_001_reset_out_reset), // reset.reset_n
		.in_ready  (fifo_0_out_ready),                    //    in.ready
		.in_valid  (fifo_0_out_valid),                    //      .valid
		.in_data   (fifo_0_out_data),                     //      .data
		.out_ready (timing_adapter_out_ready),            //   out.ready
		.out_valid (timing_adapter_out_valid),            //      .valid
		.out_data  (timing_adapter_out_data)              //      .data
	);

	demo_de0_sys_timer_0 timer_0 (
		.clk        (altpll_0_c0_clk),                                      //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                  // reset.reset_n
		.address    (timer_0_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_0_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_0_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_0_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_0_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                              //   irq.irq
	);

	demo_de0_sys_spi_0 spi_0 (
		.clk           (altpll_0_c0_clk),                                                  //              clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                              //            reset.reset_n
		.data_from_cpu (spi_0_spi_control_port_translator_avalon_anti_slave_0_writedata),  // spi_control_port.writedata
		.data_to_cpu   (spi_0_spi_control_port_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.mem_addr      (spi_0_spi_control_port_translator_avalon_anti_slave_0_address),    //                 .address
		.read_n        (~spi_0_spi_control_port_translator_avalon_anti_slave_0_read),      //                 .read_n
		.spi_select    (spi_0_spi_control_port_translator_avalon_anti_slave_0_chipselect), //                 .chipselect
		.write_n       (~spi_0_spi_control_port_translator_avalon_anti_slave_0_write),     //                 .write_n
		.dataavailable (),                                                                 //                 .dataavailable
		.endofpacket   (),                                                                 //                 .endofpacket
		.readyfordata  (),                                                                 //                 .readyfordata
		.irq           (irq_mapper_receiver3_irq),                                         //              irq.irq
		.MISO          (sdcard_MISO),                                                      //         external.export
		.MOSI          (sdcard_MOSI),                                                      //                 .export
		.SCLK          (sdcard_SCLK),                                                      //                 .export
		.SS_n          (sdcard_SS_n)                                                       //                 .export
	);

	demo_de0_sys_pio_0 pio_0 (
		.clk      (altpll_0_c0_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),              //               reset.reset_n
		.address  (pio_0_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (pio_0_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (sw_export)                                         // external_connection.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (25),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_0_instruction_master_translator (
		.clk                   (altpll_0_c0_clk),                                                                    //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                 //                     reset.reset
		.uav_address           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_qsys_0_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_qsys_0_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (nios2_qsys_0_instruction_master_read),                                               //                          .read
		.av_readdata           (nios2_qsys_0_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount         (1'b1),                                                                               //               (terminated)
		.av_byteenable         (4'b1111),                                                                            //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                                               //               (terminated)
		.av_readdatavalid      (),                                                                                   //               (terminated)
		.av_write              (1'b0),                                                                               //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                               //               (terminated)
		.av_lock               (1'b0),                                                                               //               (terminated)
		.av_debugaccess        (1'b0),                                                                               //               (terminated)
		.uav_clken             (),                                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                                //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (25),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) nios2_qsys_0_data_master_translator (
		.clk                   (altpll_0_c0_clk),                                                             //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                          //                     reset.reset
		.uav_address           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_qsys_0_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_qsys_0_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_qsys_0_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_qsys_0_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (nios2_qsys_0_data_master_byteenable),                                         //                          .byteenable
		.av_read               (nios2_qsys_0_data_master_read),                                               //                          .read
		.av_readdata           (nios2_qsys_0_data_master_readdata),                                           //                          .readdata
		.av_write              (nios2_qsys_0_data_master_write),                                              //                          .write
		.av_writedata          (nios2_qsys_0_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (nios2_qsys_0_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_readdatavalid      (),                                                                            //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_qsys_0_jtag_debug_module_translator (
		.clk                   (altpll_0_c0_clk),                                                                           //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                        //                    reset.reset
		.uav_address           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                                          //              (terminated)
		.av_burstcount         (),                                                                                          //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                      //              (terminated)
		.av_waitrequest        (1'b0),                                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                                          //              (terminated)
		.av_lock               (),                                                                                          //              (terminated)
		.av_clken              (),                                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                                      //              (terminated)
		.av_outputenable       ()                                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (11),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ram_0_s1_translator (
		.clk                   (altpll_0_c0_clk),                                                     //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                  //                    reset.reset
		.uav_address           (ram_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ram_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ram_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ram_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ram_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (ram_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ram_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (ram_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (ram_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (ram_0_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                    //              (terminated)
		.av_begintransfer      (),                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                    //              (terminated)
		.av_burstcount         (),                                                                    //              (terminated)
		.av_readdatavalid      (1'b0),                                                                //              (terminated)
		.av_waitrequest        (1'b0),                                                                //              (terminated)
		.av_writebyteenable    (),                                                                    //              (terminated)
		.av_lock               (),                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                //              (terminated)
		.av_debugaccess        (),                                                                    //              (terminated)
		.av_outputenable       ()                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (2),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (1),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) rom_0_uas_translator (
		.clk                   (altpll_0_c0_clk),                                                      //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                   //                    reset.reset
		.uav_address           (rom_0_uas_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (rom_0_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (rom_0_uas_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (rom_0_uas_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (rom_0_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (rom_0_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (rom_0_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (rom_0_uas_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (rom_0_uas_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (rom_0_uas_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (rom_0_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (rom_0_uas_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (rom_0_uas_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (rom_0_uas_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (rom_0_uas_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (rom_0_uas_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (rom_0_uas_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (rom_0_uas_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (rom_0_uas_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (rom_0_uas_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_lock               (rom_0_uas_translator_avalon_anti_slave_0_lock),                        //                         .lock
		.av_debugaccess        (rom_0_uas_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_qsys_0_control_slave_translator (
		.clk                   (altpll_0_c0_clk),                                                                       //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                    //                    reset.reset
		.uav_address           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                                      //              (terminated)
		.av_read               (),                                                                                      //              (terminated)
		.av_writedata          (),                                                                                      //              (terminated)
		.av_begintransfer      (),                                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                                      //              (terminated)
		.av_burstcount         (),                                                                                      //              (terminated)
		.av_byteenable         (),                                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                                      //              (terminated)
		.av_lock               (),                                                                                      //              (terminated)
		.av_chipselect         (),                                                                                      //              (terminated)
		.av_clken              (),                                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                                  //              (terminated)
		.av_debugaccess        (),                                                                                      //              (terminated)
		.av_outputenable       ()                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) altpll_0_pll_slave_translator (
		.clk                   (clk_clk),                                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                //                    reset.reset
		.uav_address           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (altpll_0_pll_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (altpll_0_pll_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (altpll_0_pll_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (altpll_0_pll_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (altpll_0_pll_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_waitrequest        (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_0_in_translator (
		.clk                   (altpll_0_c0_clk),                                                      //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                   //                    reset.reset
		.uav_address           (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (fifo_0_in_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (fifo_0_in_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_writedata          (fifo_0_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (fifo_0_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_read               (),                                                                     //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                 //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_0_in_csr_translator (
		.clk                   (altpll_0_c0_clk),                                                          //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address           (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (fifo_0_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (fifo_0_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (fifo_0_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (fifo_0_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (fifo_0_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) m2vdec_0_control_translator (
		.clk                   (altpll_0_c0_clk),                                                             //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                          //                    reset.reset
		.uav_address           (m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (m2vdec_0_control_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (m2vdec_0_control_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (m2vdec_0_control_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (m2vdec_0_control_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (m2vdec_0_control_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_readdatavalid      (m2vdec_0_control_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_byteenable         (),                                                                            //              (terminated)
		.av_waitrequest        (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.av_chipselect         (),                                                                            //              (terminated)
		.av_clken              (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hexdisp_0_ctrl_translator (
		.clk                   (altpll_0_c0_clk),                                                           //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                        //                    reset.reset
		.uav_address           (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (hexdisp_0_ctrl_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (hexdisp_0_ctrl_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_writedata          (hexdisp_0_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_read               (),                                                                          //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                      //              (terminated)
		.av_begintransfer      (),                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                          //              (terminated)
		.av_burstcount         (),                                                                          //              (terminated)
		.av_byteenable         (),                                                                          //              (terminated)
		.av_readdatavalid      (1'b0),                                                                      //              (terminated)
		.av_waitrequest        (1'b0),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                          //              (terminated)
		.av_lock               (),                                                                          //              (terminated)
		.av_chipselect         (),                                                                          //              (terminated)
		.av_clken              (),                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                      //              (terminated)
		.av_debugaccess        (),                                                                          //              (terminated)
		.av_outputenable       ()                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) m2vdd_hx8347a_0_ctrl_translator (
		.clk                   (altpll_0_c0_clk),                                                                 //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                              //                    reset.reset
		.uav_address           (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (m2vdd_hx8347a_0_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (m2vdd_hx8347a_0_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (m2vdd_hx8347a_0_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (m2vdd_hx8347a_0_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_readdatavalid      (m2vdd_hx8347a_0_ctrl_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (m2vdd_hx8347a_0_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                                //              (terminated)
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_byteenable         (),                                                                                //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.av_chipselect         (),                                                                                //              (terminated)
		.av_clken              (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_0_s1_translator (
		.clk                   (altpll_0_c0_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) spi_0_spi_control_port_translator (
		.clk                   (altpll_0_c0_clk),                                                                   //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                //                    reset.reset
		.uav_address           (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (spi_0_spi_control_port_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (spi_0_spi_control_port_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (spi_0_spi_control_port_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (spi_0_spi_control_port_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (spi_0_spi_control_port_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (spi_0_spi_control_port_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                  //              (terminated)
		.av_byteenable         (),                                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                                              //              (terminated)
		.av_waitrequest        (1'b0),                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                                  //              (terminated)
		.av_lock               (),                                                                                  //              (terminated)
		.av_clken              (),                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                              //              (terminated)
		.av_debugaccess        (),                                                                                  //              (terminated)
		.av_outputenable       ()                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_0_s1_translator (
		.clk                   (altpll_0_c0_clk),                                                     //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                  //                    reset.reset
		.uav_address           (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pio_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (pio_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                    //              (terminated)
		.av_read               (),                                                                    //              (terminated)
		.av_writedata          (),                                                                    //              (terminated)
		.av_begintransfer      (),                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                    //              (terminated)
		.av_burstcount         (),                                                                    //              (terminated)
		.av_byteenable         (),                                                                    //              (terminated)
		.av_readdatavalid      (1'b0),                                                                //              (terminated)
		.av_waitrequest        (1'b0),                                                                //              (terminated)
		.av_writebyteenable    (),                                                                    //              (terminated)
		.av_lock               (),                                                                    //              (terminated)
		.av_chipselect         (),                                                                    //              (terminated)
		.av_clken              (),                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                //              (terminated)
		.av_debugaccess        (),                                                                    //              (terminated)
		.av_outputenable       ()                                                                     //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (23),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (23),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) m2vdd_hx8347a_0_fbuf_translator (
		.clk                   (altpll_0_c0_clk),                                                         //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                      //                     reset.reset
		.uav_address           (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (m2vdd_hx8347a_0_fbuf_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (m2vdd_hx8347a_0_fbuf_waitrequest),                                        //                          .waitrequest
		.av_read               (m2vdd_hx8347a_0_fbuf_read),                                               //                          .read
		.av_readdata           (m2vdd_hx8347a_0_fbuf_readdata),                                           //                          .readdata
		.av_readdatavalid      (m2vdd_hx8347a_0_fbuf_readdatavalid),                                      //                          .readdatavalid
		.av_write              (m2vdd_hx8347a_0_fbuf_write),                                              //                          .write
		.av_writedata          (m2vdd_hx8347a_0_fbuf_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                    //               (terminated)
		.av_byteenable         (2'b11),                                                                   //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                    //               (terminated)
		.av_begintransfer      (1'b0),                                                                    //               (terminated)
		.av_chipselect         (1'b0),                                                                    //               (terminated)
		.av_lock               (1'b0),                                                                    //               (terminated)
		.av_debugaccess        (1'b0),                                                                    //               (terminated)
		.uav_clken             (),                                                                        //               (terminated)
		.av_clken              (1'b1)                                                                     //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (23),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (23),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) m2vdec_0_fbuf_translator (
		.clk                   (altpll_0_c0_clk),                                                  //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                               //                     reset.reset
		.uav_address           (m2vdec_0_fbuf_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (m2vdec_0_fbuf_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (m2vdec_0_fbuf_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (m2vdec_0_fbuf_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (m2vdec_0_fbuf_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (m2vdec_0_fbuf_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (m2vdec_0_fbuf_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (m2vdec_0_fbuf_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (m2vdec_0_fbuf_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (m2vdec_0_fbuf_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (m2vdec_0_fbuf_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (m2vdec_0_fbuf_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (m2vdec_0_fbuf_waitrequest),                                        //                          .waitrequest
		.av_read               (m2vdec_0_fbuf_read),                                               //                          .read
		.av_readdata           (m2vdec_0_fbuf_readdata),                                           //                          .readdata
		.av_readdatavalid      (m2vdec_0_fbuf_readdatavalid),                                      //                          .readdatavalid
		.av_write              (m2vdec_0_fbuf_write),                                              //                          .write
		.av_writedata          (m2vdec_0_fbuf_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                             //               (terminated)
		.av_byteenable         (2'b11),                                                            //               (terminated)
		.av_beginbursttransfer (1'b0),                                                             //               (terminated)
		.av_begintransfer      (1'b0),                                                             //               (terminated)
		.av_chipselect         (1'b0),                                                             //               (terminated)
		.av_lock               (1'b0),                                                             //               (terminated)
		.av_debugaccess        (1'b0),                                                             //               (terminated)
		.uav_clken             (),                                                                 //               (terminated)
		.av_clken              (1'b1)                                                              //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (23),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_0_s1_translator (
		.clk                   (altpll_0_c0_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address           (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sdram_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sdram_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sdram_0_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sdram_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sdram_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sdram_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (sdram_0_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (sdram_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (81),
		.PKT_PROTECTION_L          (81),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pio_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                               //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src12_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src12_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src12_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src12_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src12_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src12_channel),                                              //                .channel
		.rf_sink_ready           (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (54),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_POSTED          (44),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.PKT_TRANS_LOCK            (47),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (55),
		.PKT_DEST_ID_H             (62),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (53),
		.PKT_BURSTWRAP_L           (51),
		.PKT_BYTE_CNT_H            (50),
		.PKT_BYTE_CNT_L            (48),
		.PKT_PROTECTION_H          (63),
		.PKT_PROTECTION_L          (63),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (64),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) rom_0_uas_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (rom_0_uas_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (rom_0_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (rom_0_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (rom_0_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (rom_0_uas_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (rom_0_uas_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (rom_0_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (rom_0_uas_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (rom_0_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (rom_0_uas_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (rom_0_uas_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (rom_0_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (rom_0_uas_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (rom_0_uas_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (rom_0_uas_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (rom_0_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                    //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                    //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                     //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                              //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                  //                .channel
		.rf_sink_ready           (rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (rom_0_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (rom_0_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (rom_0_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (rom_0_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (rom_0_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (rom_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (rom_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (rom_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (rom_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (rom_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (rom_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (65),
		.FIFO_DEPTH          (4),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.in_data           (rom_0_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (rom_0_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (rom_0_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (rom_0_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (rom_0_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (rom_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (81),
		.PKT_PROTECTION_L          (81),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) spi_0_spi_control_port_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src11_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src11_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_001_src11_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src11_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src11_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src11_channel),                                                            //                .channel
		.rf_sink_ready           (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (81),
		.PKT_PROTECTION_L          (81),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                     //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                                     //                .channel
		.rf_sink_ready           (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                     //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (81),
		.PKT_PROTECTION_L          (81),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) m2vdec_0_control_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (m2vdec_0_control_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                                       //                .channel
		.rf_sink_ready           (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                       //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (81),
		.PKT_PROTECTION_L          (81),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src10_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src10_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src10_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src10_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src10_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src10_channel),                                                //                .channel
		.rf_sink_ready           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (81),
		.PKT_PROTECTION_L          (81),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ram_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                               //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (ram_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ram_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ram_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ram_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                  //                .channel
		.rf_sink_ready           (ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (ram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (81),
		.PKT_PROTECTION_L          (81),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) altpll_0_pll_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_out_ready),                                                                       //              cp.ready
		.cp_valid                (crosser_out_valid),                                                                       //                .valid
		.cp_data                 (crosser_out_data),                                                                        //                .data
		.cp_startofpacket        (crosser_out_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (crosser_out_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (crosser_out_channel),                                                                     //                .channel
		.rf_sink_ready           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_startofpacket  (1'b0),                                                                              // (terminated)
		.in_endofpacket    (1'b0),                                                                              // (terminated)
		.out_startofpacket (),                                                                                  // (terminated)
		.out_endofpacket   (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (81),
		.PKT_PROTECTION_L          (81),
		.PKT_BEGIN_BURST           (72),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.ST_DATA_W                 (82),
		.ST_CHANNEL_W              (13),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7)
	) nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent (
		.clk              (altpll_0_c0_clk),                                                                      //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.av_address       (nios2_qsys_0_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_001_src_valid),                                                           //        rp.valid
		.rp_data          (rsp_xbar_mux_001_src_data),                                                            //          .data
		.rp_channel       (rsp_xbar_mux_001_src_channel),                                                         //          .channel
		.rp_startofpacket (rsp_xbar_mux_001_src_startofpacket),                                                   //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_001_src_endofpacket),                                                     //          .endofpacket
		.rp_ready         (rsp_xbar_mux_001_src_ready)                                                            //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (81),
		.PKT_PROTECTION_L          (81),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_0_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                    //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                    //                .channel
		.rf_sink_ready           (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (81),
		.PKT_PROTECTION_L          (81),
		.PKT_BEGIN_BURST           (72),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.ST_DATA_W                 (82),
		.ST_CHANNEL_W              (13),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (3)
	) nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (altpll_0_c0_clk),                                                                             //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                          // clk_reset.reset
		.av_address       (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_src_valid),                                                                      //        rp.valid
		.rp_data          (rsp_xbar_mux_src_data),                                                                       //          .data
		.rp_channel       (rsp_xbar_mux_src_channel),                                                                    //          .channel
		.rp_startofpacket (rsp_xbar_mux_src_startofpacket),                                                              //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_src_endofpacket),                                                                //          .endofpacket
		.rp_ready         (rsp_xbar_mux_src_ready)                                                                       //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (81),
		.PKT_PROTECTION_L          (81),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                                                 //                .channel
		.rf_sink_ready           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (81),
		.PKT_PROTECTION_L          (81),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src9_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src9_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_001_src9_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src9_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src9_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src9_channel),                                                           //                .channel
		.rf_sink_ready           (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (81),
		.PKT_PROTECTION_L          (81),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                  //       clk_reset.reset
		.m0_address              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                              //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                              //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                               //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                            //                .channel
		.rf_sink_ready           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                  // clk_reset.reset
		.in_data           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (69),
		.PKT_BYTE_CNT_H            (68),
		.PKT_BYTE_CNT_L            (66),
		.PKT_PROTECTION_H          (81),
		.PKT_PROTECTION_L          (81),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fifo_0_in_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_0_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_0_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_0_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_0_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                //                .channel
		.rf_sink_ready           (fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_0_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.in_data           (fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_0_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_0_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (53),
		.PKT_PROTECTION_L          (53),
		.PKT_BEGIN_BURST           (50),
		.PKT_BURSTWRAP_H           (49),
		.PKT_BURSTWRAP_L           (48),
		.PKT_BYTE_CNT_H            (47),
		.PKT_BYTE_CNT_L            (46),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (51),
		.PKT_SRC_ID_L              (51),
		.PKT_DEST_ID_H             (52),
		.PKT_DEST_ID_L             (52),
		.ST_DATA_W                 (54),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (3)
	) m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent (
		.clk              (altpll_0_c0_clk),                                                                  //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.av_address       (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_013_src0_valid),                                                    //        rp.valid
		.rp_data          (rsp_xbar_demux_013_src0_data),                                                     //          .data
		.rp_channel       (rsp_xbar_demux_013_src0_channel),                                                  //          .channel
		.rp_startofpacket (rsp_xbar_demux_013_src0_startofpacket),                                            //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),                                              //          .endofpacket
		.rp_ready         (rsp_xbar_demux_013_src0_ready)                                                     //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (50),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (51),
		.PKT_SRC_ID_L              (51),
		.PKT_DEST_ID_H             (52),
		.PKT_DEST_ID_L             (52),
		.PKT_BURSTWRAP_H           (49),
		.PKT_BURSTWRAP_L           (48),
		.PKT_BYTE_CNT_H            (47),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (53),
		.PKT_PROTECTION_L          (53),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (54),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sdram_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_013_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_013_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_013_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_013_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_013_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_013_src_channel),                                                    //                .channel
		.rf_sink_ready           (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (55),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (53),
		.PKT_PROTECTION_L          (53),
		.PKT_BEGIN_BURST           (50),
		.PKT_BURSTWRAP_H           (49),
		.PKT_BURSTWRAP_L           (48),
		.PKT_BYTE_CNT_H            (47),
		.PKT_BYTE_CNT_L            (46),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (51),
		.PKT_SRC_ID_L              (51),
		.PKT_DEST_ID_H             (52),
		.PKT_DEST_ID_L             (52),
		.ST_DATA_W                 (54),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3)
	) m2vdec_0_fbuf_translator_avalon_universal_master_0_agent (
		.clk              (altpll_0_c0_clk),                                                           //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                        // clk_reset.reset
		.av_address       (m2vdec_0_fbuf_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (m2vdec_0_fbuf_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (m2vdec_0_fbuf_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (m2vdec_0_fbuf_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (m2vdec_0_fbuf_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (m2vdec_0_fbuf_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (m2vdec_0_fbuf_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (m2vdec_0_fbuf_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (m2vdec_0_fbuf_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (m2vdec_0_fbuf_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (m2vdec_0_fbuf_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (m2vdec_0_fbuf_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (m2vdec_0_fbuf_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (m2vdec_0_fbuf_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (m2vdec_0_fbuf_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (m2vdec_0_fbuf_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_013_src1_valid),                                             //        rp.valid
		.rp_data          (rsp_xbar_demux_013_src1_data),                                              //          .data
		.rp_channel       (rsp_xbar_demux_013_src1_channel),                                           //          .channel
		.rp_startofpacket (rsp_xbar_demux_013_src1_startofpacket),                                     //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_013_src1_endofpacket),                                       //          .endofpacket
		.rp_ready         (rsp_xbar_demux_013_src1_ready)                                              //          .ready
	);

	demo_de0_sys_addr_router addr_router (
		.sink_ready         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                       //       src.ready
		.src_valid          (addr_router_src_valid),                                                                       //          .valid
		.src_data           (addr_router_src_data),                                                                        //          .data
		.src_channel        (addr_router_src_channel),                                                                     //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                                  //          .endofpacket
	);

	demo_de0_sys_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                            //          .valid
		.src_data           (addr_router_001_src_data),                                                             //          .data
		.src_channel        (addr_router_001_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                       //          .endofpacket
	);

	demo_de0_sys_id_router id_router (
		.sink_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                           //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                       //       src.ready
		.src_valid          (id_router_src_valid),                                                                       //          .valid
		.src_data           (id_router_src_data),                                                                        //          .data
		.src_channel        (id_router_src_channel),                                                                     //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                                  //          .endofpacket
	);

	demo_de0_sys_id_router id_router_001 (
		.sink_ready         (ram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ram_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                             //       src.ready
		.src_valid          (id_router_001_src_valid),                                             //          .valid
		.src_data           (id_router_001_src_data),                                              //          .data
		.src_channel        (id_router_001_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                        //          .endofpacket
	);

	demo_de0_sys_id_router_002 id_router_002 (
		.sink_ready         (rom_0_uas_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (rom_0_uas_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (rom_0_uas_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (rom_0_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (rom_0_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                              //       src.ready
		.src_valid          (id_router_002_src_valid),                                              //          .valid
		.src_data           (id_router_002_src_data),                                               //          .data
		.src_channel        (id_router_002_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                         //          .endofpacket
	);

	demo_de0_sys_id_router_003 id_router_003 (
		.sink_ready         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                               //       src.ready
		.src_valid          (id_router_003_src_valid),                                                               //          .valid
		.src_data           (id_router_003_src_data),                                                                //          .data
		.src_channel        (id_router_003_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                          //          .endofpacket
	);

	demo_de0_sys_id_router_003 id_router_004 (
		.sink_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                       //       src.ready
		.src_valid          (id_router_004_src_valid),                                                       //          .valid
		.src_data           (id_router_004_src_data),                                                        //          .data
		.src_channel        (id_router_004_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                  //          .endofpacket
	);

	demo_de0_sys_id_router_003 id_router_005 (
		.sink_ready         (fifo_0_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_0_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_0_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_0_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_0_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                              //       src.ready
		.src_valid          (id_router_005_src_valid),                                              //          .valid
		.src_data           (id_router_005_src_data),                                               //          .data
		.src_channel        (id_router_005_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                         //          .endofpacket
	);

	demo_de0_sys_id_router_003 id_router_006 (
		.sink_ready         (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_0_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                  //       src.ready
		.src_valid          (id_router_006_src_valid),                                                  //          .valid
		.src_data           (id_router_006_src_data),                                                   //          .data
		.src_channel        (id_router_006_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                             //          .endofpacket
	);

	demo_de0_sys_id_router_003 id_router_007 (
		.sink_ready         (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (m2vdec_0_control_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                     //       src.ready
		.src_valid          (id_router_007_src_valid),                                                     //          .valid
		.src_data           (id_router_007_src_data),                                                      //          .data
		.src_channel        (id_router_007_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                //          .endofpacket
	);

	demo_de0_sys_id_router_003 id_router_008 (
		.sink_ready         (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hexdisp_0_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                           //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                   //       src.ready
		.src_valid          (id_router_008_src_valid),                                                   //          .valid
		.src_data           (id_router_008_src_data),                                                    //          .data
		.src_channel        (id_router_008_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                              //          .endofpacket
	);

	demo_de0_sys_id_router_003 id_router_009 (
		.sink_ready         (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (m2vdd_hx8347a_0_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                         //       src.ready
		.src_valid          (id_router_009_src_valid),                                                         //          .valid
		.src_data           (id_router_009_src_data),                                                          //          .data
		.src_channel        (id_router_009_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                    //          .endofpacket
	);

	demo_de0_sys_id_router_003 id_router_010 (
		.sink_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                               //       src.ready
		.src_valid          (id_router_010_src_valid),                                               //          .valid
		.src_data           (id_router_010_src_data),                                                //          .data
		.src_channel        (id_router_010_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                          //          .endofpacket
	);

	demo_de0_sys_id_router_003 id_router_011 (
		.sink_ready         (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                           //       src.ready
		.src_valid          (id_router_011_src_valid),                                                           //          .valid
		.src_data           (id_router_011_src_data),                                                            //          .data
		.src_channel        (id_router_011_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                                      //          .endofpacket
	);

	demo_de0_sys_id_router_003 id_router_012 (
		.sink_ready         (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                             //       src.ready
		.src_valid          (id_router_012_src_valid),                                             //          .valid
		.src_data           (id_router_012_src_data),                                              //          .data
		.src_channel        (id_router_012_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                        //          .endofpacket
	);

	demo_de0_sys_addr_router_002 addr_router_002 (
		.sink_ready         (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (m2vdd_hx8347a_0_fbuf_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                        //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                        //          .valid
		.src_data           (addr_router_002_src_data),                                                         //          .data
		.src_channel        (addr_router_002_src_channel),                                                      //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                   //          .endofpacket
	);

	demo_de0_sys_addr_router_002 addr_router_003 (
		.sink_ready         (m2vdec_0_fbuf_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (m2vdec_0_fbuf_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (m2vdec_0_fbuf_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (m2vdec_0_fbuf_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (m2vdec_0_fbuf_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                           //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                 //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                 //          .valid
		.src_data           (addr_router_003_src_data),                                                  //          .data
		.src_channel        (addr_router_003_src_channel),                                               //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                            //          .endofpacket
	);

	demo_de0_sys_id_router_013 id_router_013 (
		.sink_ready         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                               //       src.ready
		.src_valid          (id_router_013_src_valid),                                               //          .valid
		.src_data           (id_router_013_src_data),                                                //          .data
		.src_channel        (id_router_013_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                          //          .endofpacket
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (54),
		.PKT_BYTE_CNT_H            (50),
		.PKT_BYTE_CNT_L            (48),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURSTWRAP_H           (53),
		.PKT_BURSTWRAP_L           (51),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.ST_DATA_W                 (64),
		.ST_CHANNEL_W              (13),
		.OUT_BYTE_CNT_H            (49),
		.OUT_BURSTWRAP_H           (53),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (altpll_0_c0_clk),                     //       cr0.clk
		.reset                 (rst_controller_001_reset_out_reset),  // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                             // reset_in0.reset
		.reset_in1  (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                                    //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1  (~reset_reset_n),                             // reset_in1.reset
		.clk        (altpll_0_c0_clk),                            //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),         // reset_out.reset
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	demo_de0_sys_cmd_xbar_demux cmd_xbar_demux (
		.clk                (altpll_0_c0_clk),                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready         (addr_router_src_ready),              //      sink.ready
		.sink_channel       (addr_router_src_channel),            //          .channel
		.sink_data          (addr_router_src_data),               //          .data
		.sink_startofpacket (addr_router_src_startofpacket),      //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),        //          .endofpacket
		.sink_valid         (addr_router_src_valid),              //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),          //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),           //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),    //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),          //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),          //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),           //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),        //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),    //          .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),          //      src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),          //          .valid
		.src2_data          (cmd_xbar_demux_src2_data),           //          .data
		.src2_channel       (cmd_xbar_demux_src2_channel),        //          .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket)     //          .endofpacket
	);

	demo_de0_sys_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (altpll_0_c0_clk),                        //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),     // clk_reset.reset
		.sink_ready          (addr_router_001_src_ready),              //      sink.ready
		.sink_channel        (addr_router_001_src_channel),            //          .channel
		.sink_data           (addr_router_001_src_data),               //          .data
		.sink_startofpacket  (addr_router_001_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_001_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_001_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket)    //          .endofpacket
	);

	demo_de0_sys_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (altpll_0_c0_clk),                       //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	demo_de0_sys_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (altpll_0_c0_clk),                       //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	demo_de0_sys_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (altpll_0_c0_clk),                       //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	demo_de0_sys_rsp_xbar_demux rsp_xbar_demux (
		.clk                (altpll_0_c0_clk),                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready         (id_router_src_ready),                //      sink.ready
		.sink_channel       (id_router_src_channel),              //          .channel
		.sink_data          (id_router_src_data),                 //          .data
		.sink_startofpacket (id_router_src_startofpacket),        //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),          //          .endofpacket
		.sink_valid         (id_router_src_valid),                //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),          //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),           //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),    //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),          //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),          //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),           //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),        //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)     //          .endofpacket
	);

	demo_de0_sys_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	demo_de0_sys_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	demo_de0_sys_rsp_xbar_demux_003 rsp_xbar_demux_003 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	demo_de0_sys_rsp_xbar_demux_003 rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	demo_de0_sys_rsp_xbar_demux_003 rsp_xbar_demux_005 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	demo_de0_sys_rsp_xbar_demux_003 rsp_xbar_demux_006 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	demo_de0_sys_rsp_xbar_demux_003 rsp_xbar_demux_007 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	demo_de0_sys_rsp_xbar_demux_003 rsp_xbar_demux_008 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	demo_de0_sys_rsp_xbar_demux_003 rsp_xbar_demux_009 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	demo_de0_sys_rsp_xbar_demux_003 rsp_xbar_demux_010 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	demo_de0_sys_rsp_xbar_demux_003 rsp_xbar_demux_011 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	demo_de0_sys_rsp_xbar_demux_003 rsp_xbar_demux_012 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	demo_de0_sys_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (altpll_0_c0_clk),                       //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	demo_de0_sys_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (altpll_0_c0_clk),                       //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (crosser_001_out_ready),                 //     sink4.ready
		.sink4_valid          (crosser_001_out_valid),                 //          .valid
		.sink4_channel        (crosser_001_out_channel),               //          .channel
		.sink4_data           (crosser_001_out_data),                  //          .data
		.sink4_startofpacket  (crosser_001_out_startofpacket),         //          .startofpacket
		.sink4_endofpacket    (crosser_001_out_endofpacket),           //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	demo_de0_sys_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	demo_de0_sys_cmd_xbar_demux_002 cmd_xbar_demux_003 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_003_src_ready),             //      sink.ready
		.sink_channel       (addr_router_003_src_channel),           //          .channel
		.sink_data          (addr_router_003_src_data),              //          .data
		.sink_startofpacket (addr_router_003_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_003_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_003_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	demo_de0_sys_cmd_xbar_mux_013 cmd_xbar_mux_013 (
		.clk                 (altpll_0_c0_clk),                       //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_013_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_013_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_013_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_013_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_013_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_013_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_002_src0_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_003_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	demo_de0_sys_rsp_xbar_demux_013 rsp_xbar_demux_013 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_013_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_013_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_013_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_013_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_013_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_013_src1_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (68),
		.IN_PKT_BYTE_CNT_L             (66),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (71),
		.IN_PKT_BURSTWRAP_L            (69),
		.IN_ST_DATA_W                  (82),
		.OUT_PKT_ADDR_H                (42),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (50),
		.OUT_PKT_BYTE_CNT_L            (48),
		.OUT_PKT_TRANS_COMPRESSED_READ (43),
		.OUT_ST_DATA_W                 (64),
		.ST_CHANNEL_W                  (13),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk               (altpll_0_c0_clk),                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset), // clk_reset.reset
		.in_valid          (cmd_xbar_mux_002_src_valid),         //      sink.valid
		.in_channel        (cmd_xbar_mux_002_src_channel),       //          .channel
		.in_startofpacket  (cmd_xbar_mux_002_src_startofpacket), //          .startofpacket
		.in_endofpacket    (cmd_xbar_mux_002_src_endofpacket),   //          .endofpacket
		.in_ready          (cmd_xbar_mux_002_src_ready),         //          .ready
		.in_data           (cmd_xbar_mux_002_src_data),          //          .data
		.out_endofpacket   (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data          (width_adapter_src_data),             //          .data
		.out_channel       (width_adapter_src_channel),          //          .channel
		.out_valid         (width_adapter_src_valid),            //          .valid
		.out_ready         (width_adapter_src_ready),            //          .ready
		.out_startofpacket (width_adapter_src_startofpacket)     //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (42),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (50),
		.IN_PKT_BYTE_CNT_L             (48),
		.IN_PKT_TRANS_COMPRESSED_READ  (43),
		.IN_PKT_BURSTWRAP_H            (53),
		.IN_PKT_BURSTWRAP_L            (51),
		.IN_ST_DATA_W                  (64),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (68),
		.OUT_PKT_BYTE_CNT_L            (66),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_ST_DATA_W                 (82),
		.ST_CHANNEL_W                  (13),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_001 (
		.clk               (altpll_0_c0_clk),                     //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),  // clk_reset.reset
		.in_valid          (id_router_002_src_valid),             //      sink.valid
		.in_channel        (id_router_002_src_channel),           //          .channel
		.in_startofpacket  (id_router_002_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_002_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_002_src_ready),             //          .ready
		.in_data           (id_router_002_src_data),              //          .data
		.out_endofpacket   (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_001_src_data),          //          .data
		.out_channel       (width_adapter_001_src_channel),       //          .channel
		.out_valid         (width_adapter_001_src_valid),         //          .valid
		.out_ready         (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket (width_adapter_001_src_startofpacket)  //          .startofpacket
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (82),
		.BITS_PER_SYMBOL     (82),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (13),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (altpll_0_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src4_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src4_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src4_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src4_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src4_data),          //              .data
		.out_ready         (crosser_out_ready),                     //           out.ready
		.out_valid         (crosser_out_valid),                     //              .valid
		.out_startofpacket (crosser_out_startofpacket),             //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),               //              .endofpacket
		.out_channel       (crosser_out_channel),                   //              .channel
		.out_data          (crosser_out_data),                      //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (82),
		.BITS_PER_SYMBOL     (82),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (13),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (altpll_0_c0_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_004_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_004_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_004_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_004_src0_data),          //              .data
		.out_ready         (crosser_001_out_ready),                 //           out.ready
		.out_valid         (crosser_001_out_valid),                 //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_001_out_channel),               //              .channel
		.out_data          (crosser_001_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	demo_de0_sys_irq_mapper irq_mapper (
		.clk           (altpll_0_c0_clk),                    //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)              //    sender.irq
	);

endmodule
